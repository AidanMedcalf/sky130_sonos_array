magic
tech sky130A
timestamp 1686033482
<< error_p >>
rect -80 77037 3274 77140
rect -80 77031 63 77037
rect -80 76987 117 77031
rect 171 76987 261 77031
rect 315 76987 405 77031
rect 459 76987 549 77031
rect 603 76987 693 77031
rect 747 76987 837 77031
rect 891 76987 981 77031
rect 1035 76987 1125 77031
rect 1252 76987 1342 77031
rect 1396 76987 1486 77031
rect 1540 76987 1630 77031
rect 1684 76987 1774 77031
rect 1828 76987 1918 77031
rect 1972 76987 2062 77031
rect 2116 76987 2206 77031
rect 2260 76987 2350 77031
rect 2477 76987 2567 77031
rect 2621 76987 2711 77031
rect 2765 76987 2855 77031
rect 2909 76987 2999 77031
rect 3053 76987 3143 77031
rect 3197 76987 3274 77031
rect -80 76793 63 76987
rect -80 76749 117 76793
rect 171 76749 261 76793
rect 315 76749 405 76793
rect 459 76749 549 76793
rect 603 76749 693 76793
rect 747 76749 837 76793
rect 891 76749 981 76793
rect 1035 76749 1125 76793
rect 1252 76749 1342 76793
rect 1396 76749 1486 76793
rect 1540 76749 1630 76793
rect 1684 76749 1774 76793
rect 1828 76749 1918 76793
rect 1972 76749 2062 76793
rect 2116 76749 2206 76793
rect 2260 76749 2350 76793
rect 2477 76749 2567 76793
rect 2621 76749 2711 76793
rect 2765 76749 2855 76793
rect 2909 76749 2999 76793
rect 3053 76749 3143 76793
rect 3197 76749 3274 76793
rect -80 76685 63 76749
rect -80 76641 117 76685
rect 171 76641 261 76685
rect 315 76641 405 76685
rect 459 76641 549 76685
rect 603 76641 693 76685
rect 747 76641 837 76685
rect 891 76641 981 76685
rect 1035 76641 1125 76685
rect 1252 76641 1342 76685
rect 1396 76641 1486 76685
rect 1540 76641 1630 76685
rect 1684 76641 1774 76685
rect 1828 76641 1918 76685
rect 1972 76641 2062 76685
rect 2116 76641 2206 76685
rect 2260 76641 2350 76685
rect 2477 76641 2567 76685
rect 2621 76641 2711 76685
rect 2765 76641 2855 76685
rect 2909 76641 2999 76685
rect 3053 76641 3143 76685
rect 3197 76641 3274 76685
rect -80 76447 63 76641
rect -80 76403 117 76447
rect 171 76403 261 76447
rect 315 76403 405 76447
rect 459 76403 549 76447
rect 603 76403 693 76447
rect 747 76403 837 76447
rect 891 76403 981 76447
rect 1035 76403 1125 76447
rect 1252 76403 1342 76447
rect 1396 76403 1486 76447
rect 1540 76403 1630 76447
rect 1684 76403 1774 76447
rect 1828 76403 1918 76447
rect 1972 76403 2062 76447
rect 2116 76403 2206 76447
rect 2260 76403 2350 76447
rect 2477 76403 2567 76447
rect 2621 76403 2711 76447
rect 2765 76403 2855 76447
rect 2909 76403 2999 76447
rect 3053 76403 3143 76447
rect 3197 76403 3274 76447
rect -80 76339 63 76403
rect -80 76295 117 76339
rect 171 76295 261 76339
rect 315 76295 405 76339
rect 459 76295 549 76339
rect 603 76295 693 76339
rect 747 76295 837 76339
rect 891 76295 981 76339
rect 1035 76295 1125 76339
rect 1252 76295 1342 76339
rect 1396 76295 1486 76339
rect 1540 76295 1630 76339
rect 1684 76295 1774 76339
rect 1828 76295 1918 76339
rect 1972 76295 2062 76339
rect 2116 76295 2206 76339
rect 2260 76295 2350 76339
rect 2477 76295 2567 76339
rect 2621 76295 2711 76339
rect 2765 76295 2855 76339
rect 2909 76295 2999 76339
rect 3053 76295 3143 76339
rect 3197 76295 3274 76339
rect -80 76101 63 76295
rect -80 76057 117 76101
rect 171 76057 261 76101
rect 315 76057 405 76101
rect 459 76057 549 76101
rect 603 76057 693 76101
rect 747 76057 837 76101
rect 891 76057 981 76101
rect 1035 76057 1125 76101
rect 1252 76057 1342 76101
rect 1396 76057 1486 76101
rect 1540 76057 1630 76101
rect 1684 76057 1774 76101
rect 1828 76057 1918 76101
rect 1972 76057 2062 76101
rect 2116 76057 2206 76101
rect 2260 76057 2350 76101
rect 2477 76057 2567 76101
rect 2621 76057 2711 76101
rect 2765 76057 2855 76101
rect 2909 76057 2999 76101
rect 3053 76057 3143 76101
rect 3197 76057 3274 76101
rect -80 75993 63 76057
rect -80 75949 117 75993
rect 171 75949 261 75993
rect 315 75949 405 75993
rect 459 75949 549 75993
rect 603 75949 693 75993
rect 747 75949 837 75993
rect 891 75949 981 75993
rect 1035 75949 1125 75993
rect 1252 75949 1342 75993
rect 1396 75949 1486 75993
rect 1540 75949 1630 75993
rect 1684 75949 1774 75993
rect 1828 75949 1918 75993
rect 1972 75949 2062 75993
rect 2116 75949 2206 75993
rect 2260 75949 2350 75993
rect 2477 75949 2567 75993
rect 2621 75949 2711 75993
rect 2765 75949 2855 75993
rect 2909 75949 2999 75993
rect 3053 75949 3143 75993
rect 3197 75949 3274 75993
rect -80 75755 63 75949
rect -80 75711 117 75755
rect 171 75711 261 75755
rect 315 75711 405 75755
rect 459 75711 549 75755
rect 603 75711 693 75755
rect 747 75711 837 75755
rect 891 75711 981 75755
rect 1035 75711 1125 75755
rect 1252 75711 1342 75755
rect 1396 75711 1486 75755
rect 1540 75711 1630 75755
rect 1684 75711 1774 75755
rect 1828 75711 1918 75755
rect 1972 75711 2062 75755
rect 2116 75711 2206 75755
rect 2260 75711 2350 75755
rect 2477 75711 2567 75755
rect 2621 75711 2711 75755
rect 2765 75711 2855 75755
rect 2909 75711 2999 75755
rect 3053 75711 3143 75755
rect 3197 75711 3274 75755
rect -80 75518 63 75711
rect -80 75474 117 75518
rect 171 75474 261 75518
rect 315 75474 405 75518
rect 459 75474 549 75518
rect 603 75474 693 75518
rect 747 75474 837 75518
rect 891 75474 981 75518
rect 1035 75474 1125 75518
rect 1252 75474 1342 75518
rect 1396 75474 1486 75518
rect 1540 75474 1630 75518
rect 1684 75474 1774 75518
rect 1828 75474 1918 75518
rect 1972 75474 2062 75518
rect 2116 75474 2206 75518
rect 2260 75474 2350 75518
rect 2477 75474 2567 75518
rect 2621 75474 2711 75518
rect 2765 75474 2855 75518
rect 2909 75474 2999 75518
rect 3053 75474 3143 75518
rect 3197 75474 3274 75518
rect -80 75280 63 75474
rect -80 75236 117 75280
rect 171 75236 261 75280
rect 315 75236 405 75280
rect 459 75236 549 75280
rect 603 75236 693 75280
rect 747 75236 837 75280
rect 891 75236 981 75280
rect 1035 75236 1125 75280
rect 1252 75236 1342 75280
rect 1396 75236 1486 75280
rect 1540 75236 1630 75280
rect 1684 75236 1774 75280
rect 1828 75236 1918 75280
rect 1972 75236 2062 75280
rect 2116 75236 2206 75280
rect 2260 75236 2350 75280
rect 2477 75236 2567 75280
rect 2621 75236 2711 75280
rect 2765 75236 2855 75280
rect 2909 75236 2999 75280
rect 3053 75236 3143 75280
rect 3197 75236 3274 75280
rect -80 75174 63 75236
rect -40 3433 117 3456
rect 171 3433 261 3456
rect 315 3433 405 3456
rect 459 3433 549 3456
rect 603 3433 693 3456
rect 747 3433 837 3456
rect 891 3433 981 3456
rect 1035 3433 1125 3456
rect 1252 3433 1342 3456
rect 1396 3433 1486 3456
rect 1540 3433 1630 3456
rect 1684 3433 1774 3456
rect 1828 3433 1918 3456
rect 1972 3433 2062 3456
rect 2116 3433 2206 3456
rect 2260 3433 2350 3456
rect 2477 3433 2567 3456
rect 2621 3433 2711 3456
rect 2765 3433 2855 3456
rect 2909 3433 2999 3456
rect 3053 3433 3143 3456
rect 3197 3433 3274 3456
rect 60628 3433 60718 3456
rect 60772 3433 60862 3456
rect 60916 3433 61006 3456
rect 61060 3433 61150 3456
rect 61277 3433 61367 3456
rect 61421 3433 61511 3456
rect 61565 3433 61655 3456
rect 61709 3433 61799 3456
rect 61853 3433 61943 3456
rect 61997 3433 62087 3456
rect 62141 3433 62231 3456
rect 62285 3433 62500 3456
rect -40 3369 63 3433
rect 62357 3369 62500 3433
rect -40 3325 117 3369
rect 171 3325 261 3369
rect 315 3325 405 3369
rect 459 3325 549 3369
rect 603 3325 693 3369
rect 747 3325 837 3369
rect 891 3325 981 3369
rect 1035 3325 1125 3369
rect 1252 3325 1342 3369
rect 1396 3325 1486 3369
rect 1540 3325 1630 3369
rect 1684 3325 1774 3369
rect 1828 3325 1918 3369
rect 1972 3325 2062 3369
rect 2116 3325 2206 3369
rect 2260 3325 2350 3369
rect 2477 3325 2567 3369
rect 2621 3325 2711 3369
rect 2765 3325 2855 3369
rect 2909 3325 2999 3369
rect 3053 3325 3143 3369
rect 3197 3325 3274 3369
rect 60628 3325 60718 3369
rect 60772 3325 60862 3369
rect 60916 3325 61006 3369
rect 61060 3325 61150 3369
rect 61277 3325 61367 3369
rect 61421 3325 61511 3369
rect 61565 3325 61655 3369
rect 61709 3325 61799 3369
rect 61853 3325 61943 3369
rect 61997 3325 62087 3369
rect 62141 3325 62231 3369
rect 62285 3325 62500 3369
rect -40 3131 63 3325
rect 62357 3131 62500 3325
rect -40 3087 117 3131
rect 171 3087 261 3131
rect 315 3087 405 3131
rect 459 3087 549 3131
rect 603 3087 693 3131
rect 747 3087 837 3131
rect 891 3087 981 3131
rect 1035 3087 1125 3131
rect 1252 3087 1342 3131
rect 1396 3087 1486 3131
rect 1540 3087 1630 3131
rect 1684 3087 1774 3131
rect 1828 3087 1918 3131
rect 1972 3087 2062 3131
rect 2116 3087 2206 3131
rect 2260 3087 2350 3131
rect 2477 3087 2567 3131
rect 2621 3087 2711 3131
rect 2765 3087 2855 3131
rect 2909 3087 2999 3131
rect 3053 3087 3143 3131
rect 3197 3087 3274 3131
rect 60628 3087 60718 3131
rect 60772 3087 60862 3131
rect 60916 3087 61006 3131
rect 61060 3087 61150 3131
rect 61277 3087 61367 3131
rect 61421 3087 61511 3131
rect 61565 3087 61655 3131
rect 61709 3087 61799 3131
rect 61853 3087 61943 3131
rect 61997 3087 62087 3131
rect 62141 3087 62231 3131
rect 62285 3087 62500 3131
rect -40 2894 63 3087
rect 62357 2894 62500 3087
rect -40 2850 117 2894
rect 171 2850 261 2894
rect 315 2850 405 2894
rect 459 2850 549 2894
rect 603 2850 693 2894
rect 747 2850 837 2894
rect 891 2850 981 2894
rect 1035 2850 1125 2894
rect 1252 2850 1342 2894
rect 1396 2850 1486 2894
rect 1540 2850 1630 2894
rect 1684 2850 1774 2894
rect 1828 2850 1918 2894
rect 1972 2850 2062 2894
rect 2116 2850 2206 2894
rect 2260 2850 2350 2894
rect 2477 2850 2567 2894
rect 2621 2850 2711 2894
rect 2765 2850 2855 2894
rect 2909 2850 2999 2894
rect 3053 2850 3143 2894
rect 3197 2850 3274 2894
rect 60628 2850 60718 2894
rect 60772 2850 60862 2894
rect 60916 2850 61006 2894
rect 61060 2850 61150 2894
rect 61277 2850 61367 2894
rect 61421 2850 61511 2894
rect 61565 2850 61655 2894
rect 61709 2850 61799 2894
rect 61853 2850 61943 2894
rect 61997 2850 62087 2894
rect 62141 2850 62231 2894
rect 62285 2850 62500 2894
rect -40 2656 63 2850
rect 62357 2656 62500 2850
rect -40 2612 117 2656
rect 171 2612 261 2656
rect 315 2612 405 2656
rect 459 2612 549 2656
rect 603 2612 693 2656
rect 747 2612 837 2656
rect 891 2612 981 2656
rect 1035 2612 1125 2656
rect 1252 2612 1342 2656
rect 1396 2612 1486 2656
rect 1540 2612 1630 2656
rect 1684 2612 1774 2656
rect 1828 2612 1918 2656
rect 1972 2612 2062 2656
rect 2116 2612 2206 2656
rect 2260 2612 2350 2656
rect 2477 2612 2567 2656
rect 2621 2612 2711 2656
rect 2765 2612 2855 2656
rect 2909 2612 2999 2656
rect 3053 2612 3143 2656
rect 3197 2612 3274 2656
rect 60628 2612 60718 2656
rect 60772 2612 60862 2656
rect 60916 2612 61006 2656
rect 61060 2612 61150 2656
rect 61277 2612 61367 2656
rect 61421 2612 61511 2656
rect 61565 2612 61655 2656
rect 61709 2612 61799 2656
rect 61853 2612 61943 2656
rect 61997 2612 62087 2656
rect 62141 2612 62231 2656
rect 62285 2612 62500 2656
rect -40 2548 63 2612
rect 62357 2548 62500 2612
rect -40 2504 117 2548
rect 171 2504 261 2548
rect 315 2504 405 2548
rect 459 2504 549 2548
rect 603 2504 693 2548
rect 747 2504 837 2548
rect 891 2504 981 2548
rect 1035 2504 1125 2548
rect 1252 2504 1342 2548
rect 1396 2504 1486 2548
rect 1540 2504 1630 2548
rect 1684 2504 1774 2548
rect 1828 2504 1918 2548
rect 1972 2504 2062 2548
rect 2116 2504 2206 2548
rect 2260 2504 2350 2548
rect 2477 2504 2567 2548
rect 2621 2504 2711 2548
rect 2765 2504 2855 2548
rect 2909 2504 2999 2548
rect 3053 2504 3143 2548
rect 3197 2504 3274 2548
rect 60628 2504 60718 2548
rect 60772 2504 60862 2548
rect 60916 2504 61006 2548
rect 61060 2504 61150 2548
rect 61277 2504 61367 2548
rect 61421 2504 61511 2548
rect 61565 2504 61655 2548
rect 61709 2504 61799 2548
rect 61853 2504 61943 2548
rect 61997 2504 62087 2548
rect 62141 2504 62231 2548
rect 62285 2504 62500 2548
rect -40 2310 63 2504
rect 62357 2310 62500 2504
rect -40 2266 117 2310
rect 171 2266 261 2310
rect 315 2266 405 2310
rect 459 2266 549 2310
rect 603 2266 693 2310
rect 747 2266 837 2310
rect 891 2266 981 2310
rect 1035 2266 1125 2310
rect 1252 2266 1342 2310
rect 1396 2266 1486 2310
rect 1540 2266 1630 2310
rect 1684 2266 1774 2310
rect 1828 2266 1918 2310
rect 1972 2266 2062 2310
rect 2116 2266 2206 2310
rect 2260 2266 2350 2310
rect 2477 2266 2567 2310
rect 2621 2266 2711 2310
rect 2765 2266 2855 2310
rect 2909 2266 2999 2310
rect 3053 2266 3143 2310
rect 3197 2266 3274 2310
rect 60628 2266 60718 2310
rect 60772 2266 60862 2310
rect 60916 2266 61006 2310
rect 61060 2266 61150 2310
rect 61277 2266 61367 2310
rect 61421 2266 61511 2310
rect 61565 2266 61655 2310
rect 61709 2266 61799 2310
rect 61853 2266 61943 2310
rect 61997 2266 62087 2310
rect 62141 2266 62231 2310
rect 62285 2266 62500 2310
rect -40 2202 63 2266
rect 62357 2202 62500 2266
rect -40 2158 117 2202
rect 171 2158 261 2202
rect 315 2158 405 2202
rect 459 2158 549 2202
rect 603 2158 693 2202
rect 747 2158 837 2202
rect 891 2158 981 2202
rect 1035 2158 1125 2202
rect 1252 2158 1342 2202
rect 1396 2158 1486 2202
rect 1540 2158 1630 2202
rect 1684 2158 1774 2202
rect 1828 2158 1918 2202
rect 1972 2158 2062 2202
rect 2116 2158 2206 2202
rect 2260 2158 2350 2202
rect 2477 2158 2567 2202
rect 2621 2158 2711 2202
rect 2765 2158 2855 2202
rect 2909 2158 2999 2202
rect 3053 2158 3143 2202
rect 3197 2158 3274 2202
rect 60628 2158 60718 2202
rect 60772 2158 60862 2202
rect 60916 2158 61006 2202
rect 61060 2158 61150 2202
rect 61277 2158 61367 2202
rect 61421 2158 61511 2202
rect 61565 2158 61655 2202
rect 61709 2158 61799 2202
rect 61853 2158 61943 2202
rect 61997 2158 62087 2202
rect 62141 2158 62231 2202
rect 62285 2158 62500 2202
rect -40 1964 63 2158
rect 62357 1964 62500 2158
rect -40 1920 117 1964
rect 171 1920 261 1964
rect 315 1920 405 1964
rect 459 1920 549 1964
rect 603 1920 693 1964
rect 747 1920 837 1964
rect 891 1920 981 1964
rect 1035 1920 1125 1964
rect 1252 1920 1342 1964
rect 1396 1920 1486 1964
rect 1540 1920 1630 1964
rect 1684 1920 1774 1964
rect 1828 1920 1918 1964
rect 1972 1920 2062 1964
rect 2116 1920 2206 1964
rect 2260 1920 2350 1964
rect 2477 1920 2567 1964
rect 2621 1920 2711 1964
rect 2765 1920 2855 1964
rect 2909 1920 2999 1964
rect 3053 1920 3143 1964
rect 3197 1920 3274 1964
rect 60628 1920 60718 1964
rect 60772 1920 60862 1964
rect 60916 1920 61006 1964
rect 61060 1920 61150 1964
rect 61277 1920 61367 1964
rect 61421 1920 61511 1964
rect 61565 1920 61655 1964
rect 61709 1920 61799 1964
rect 61853 1920 61943 1964
rect 61997 1920 62087 1964
rect 62141 1920 62231 1964
rect 62285 1920 62500 1964
rect -40 1856 63 1920
rect 62357 1856 62500 1920
rect -40 1812 117 1856
rect 171 1812 261 1856
rect 315 1812 405 1856
rect 459 1812 549 1856
rect 603 1812 693 1856
rect 747 1812 837 1856
rect 891 1812 981 1856
rect 1035 1812 1125 1856
rect 1252 1812 1342 1856
rect 1396 1812 1486 1856
rect 1540 1812 1630 1856
rect 1684 1812 1774 1856
rect 1828 1812 1918 1856
rect 1972 1812 2062 1856
rect 2116 1812 2206 1856
rect 2260 1812 2350 1856
rect 2477 1812 2567 1856
rect 2621 1812 2711 1856
rect 2765 1812 2855 1856
rect 2909 1812 2999 1856
rect 3053 1812 3143 1856
rect 3197 1812 3274 1856
rect 60628 1812 60718 1856
rect 60772 1812 60862 1856
rect 60916 1812 61006 1856
rect 61060 1812 61150 1856
rect 61277 1812 61367 1856
rect 61421 1812 61511 1856
rect 61565 1812 61655 1856
rect 61709 1812 61799 1856
rect 61853 1812 61943 1856
rect 61997 1812 62087 1856
rect 62141 1812 62231 1856
rect 62285 1812 62500 1856
rect -40 1618 63 1812
rect 62357 1618 62500 1812
rect -40 1574 117 1618
rect 171 1574 261 1618
rect 315 1574 405 1618
rect 459 1574 549 1618
rect 603 1574 693 1618
rect 747 1574 837 1618
rect 891 1574 981 1618
rect 1035 1574 1125 1618
rect 1252 1574 1342 1618
rect 1396 1574 1486 1618
rect 1540 1574 1630 1618
rect 1684 1574 1774 1618
rect 1828 1574 1918 1618
rect 1972 1574 2062 1618
rect 2116 1574 2206 1618
rect 2260 1574 2350 1618
rect 2477 1574 2567 1618
rect 2621 1574 2711 1618
rect 2765 1574 2855 1618
rect 2909 1574 2999 1618
rect 3053 1574 3143 1618
rect 3197 1574 3274 1618
rect 60628 1574 60718 1618
rect 60772 1574 60862 1618
rect 60916 1574 61006 1618
rect 61060 1574 61150 1618
rect 61277 1574 61367 1618
rect 61421 1574 61511 1618
rect 61565 1574 61655 1618
rect 61709 1574 61799 1618
rect 61853 1574 61943 1618
rect 61997 1574 62087 1618
rect 62141 1574 62231 1618
rect 62285 1574 62500 1618
rect -40 1381 63 1574
rect 62357 1381 62500 1574
rect -40 1337 117 1381
rect 171 1337 261 1381
rect 315 1337 405 1381
rect 459 1337 549 1381
rect 603 1337 693 1381
rect 747 1337 837 1381
rect 891 1337 981 1381
rect 1035 1337 1125 1381
rect 1252 1337 1342 1381
rect 1396 1337 1486 1381
rect 1540 1337 1630 1381
rect 1684 1337 1774 1381
rect 1828 1337 1918 1381
rect 1972 1337 2062 1381
rect 2116 1337 2206 1381
rect 2260 1337 2350 1381
rect 2477 1337 2567 1381
rect 2621 1337 2711 1381
rect 2765 1337 2855 1381
rect 2909 1337 2999 1381
rect 3053 1337 3143 1381
rect 3197 1337 3274 1381
rect 60628 1337 60718 1381
rect 60772 1337 60862 1381
rect 60916 1337 61006 1381
rect 61060 1337 61150 1381
rect 61277 1337 61367 1381
rect 61421 1337 61511 1381
rect 61565 1337 61655 1381
rect 61709 1337 61799 1381
rect 61853 1337 61943 1381
rect 61997 1337 62087 1381
rect 62141 1337 62231 1381
rect 62285 1337 62500 1381
rect -40 1143 63 1337
rect 62357 1143 62500 1337
rect -40 1099 117 1143
rect 171 1099 261 1143
rect 315 1099 405 1143
rect 459 1099 549 1143
rect 603 1099 693 1143
rect 747 1099 837 1143
rect 891 1099 981 1143
rect 1035 1099 1125 1143
rect 1252 1099 1342 1143
rect 1396 1099 1486 1143
rect 1540 1099 1630 1143
rect 1684 1099 1774 1143
rect 1828 1099 1918 1143
rect 1972 1099 2062 1143
rect 2116 1099 2206 1143
rect 2260 1099 2350 1143
rect 2477 1099 2567 1143
rect 2621 1099 2711 1143
rect 2765 1099 2855 1143
rect 2909 1099 2999 1143
rect 3053 1099 3143 1143
rect 3197 1099 3274 1143
rect 60628 1099 60718 1143
rect 60772 1099 60862 1143
rect 60916 1099 61006 1143
rect 61060 1099 61150 1143
rect 61277 1099 61367 1143
rect 61421 1099 61511 1143
rect 61565 1099 61655 1143
rect 61709 1099 61799 1143
rect 61853 1099 61943 1143
rect 61997 1099 62087 1143
rect 62141 1099 62231 1143
rect 62285 1099 62500 1143
rect -40 1035 63 1099
rect 62357 1035 62500 1099
rect -40 991 117 1035
rect 171 991 261 1035
rect 315 991 405 1035
rect 459 991 549 1035
rect 603 991 693 1035
rect 747 991 837 1035
rect 891 991 981 1035
rect 1035 991 1125 1035
rect 1252 991 1342 1035
rect 1396 991 1486 1035
rect 1540 991 1630 1035
rect 1684 991 1774 1035
rect 1828 991 1918 1035
rect 1972 991 2062 1035
rect 2116 991 2206 1035
rect 2260 991 2350 1035
rect 2477 991 2567 1035
rect 2621 991 2711 1035
rect 2765 991 2855 1035
rect 2909 991 2999 1035
rect 3053 991 3143 1035
rect 3197 991 3274 1035
rect 60628 991 60718 1035
rect 60772 991 60862 1035
rect 60916 991 61006 1035
rect 61060 991 61150 1035
rect 61277 991 61367 1035
rect 61421 991 61511 1035
rect 61565 991 61655 1035
rect 61709 991 61799 1035
rect 61853 991 61943 1035
rect 61997 991 62087 1035
rect 62141 991 62231 1035
rect 62285 991 62500 1035
rect -40 797 63 991
rect 62357 797 62500 991
rect -40 753 117 797
rect 171 753 261 797
rect 315 753 405 797
rect 459 753 549 797
rect 603 753 693 797
rect 747 753 837 797
rect 891 753 981 797
rect 1035 753 1125 797
rect 1252 753 1342 797
rect 1396 753 1486 797
rect 1540 753 1630 797
rect 1684 753 1774 797
rect 1828 753 1918 797
rect 1972 753 2062 797
rect 2116 753 2206 797
rect 2260 753 2350 797
rect 2477 753 2567 797
rect 2621 753 2711 797
rect 2765 753 2855 797
rect 2909 753 2999 797
rect 3053 753 3143 797
rect 3197 753 3274 797
rect 60628 753 60718 797
rect 60772 753 60862 797
rect 60916 753 61006 797
rect 61060 753 61150 797
rect 61277 753 61367 797
rect 61421 753 61511 797
rect 61565 753 61655 797
rect 61709 753 61799 797
rect 61853 753 61943 797
rect 61997 753 62087 797
rect 62141 753 62231 797
rect 62285 753 62500 797
rect -40 689 63 753
rect 62357 689 62500 753
rect -40 645 117 689
rect 171 645 261 689
rect 315 645 405 689
rect 459 645 549 689
rect 603 645 693 689
rect 747 645 837 689
rect 891 645 981 689
rect 1035 645 1125 689
rect 1252 645 1342 689
rect 1396 645 1486 689
rect 1540 645 1630 689
rect 1684 645 1774 689
rect 1828 645 1918 689
rect 1972 645 2062 689
rect 2116 645 2206 689
rect 2260 645 2350 689
rect 2477 645 2567 689
rect 2621 645 2711 689
rect 2765 645 2855 689
rect 2909 645 2999 689
rect 3053 645 3143 689
rect 3197 645 3274 689
rect 60628 645 60718 689
rect 60772 645 60862 689
rect 60916 645 61006 689
rect 61060 645 61150 689
rect 61277 645 61367 689
rect 61421 645 61511 689
rect 61565 645 61655 689
rect 61709 645 61799 689
rect 61853 645 61943 689
rect 61997 645 62087 689
rect 62141 645 62231 689
rect 62285 645 62500 689
rect -40 451 63 645
rect 62357 451 62500 645
rect -40 407 117 451
rect 171 407 261 451
rect 315 407 405 451
rect 459 407 549 451
rect 603 407 693 451
rect 747 407 837 451
rect 891 407 981 451
rect 1035 407 1125 451
rect 1252 407 1342 451
rect 1396 407 1486 451
rect 1540 407 1630 451
rect 1684 407 1774 451
rect 1828 407 1918 451
rect 1972 407 2062 451
rect 2116 407 2206 451
rect 2260 407 2350 451
rect 2477 407 2567 451
rect 2621 407 2711 451
rect 2765 407 2855 451
rect 2909 407 2999 451
rect 3053 407 3143 451
rect 3197 407 3274 451
rect 60628 407 60718 451
rect 60772 407 60862 451
rect 60916 407 61006 451
rect 61060 407 61150 451
rect 61277 407 61367 451
rect 61421 407 61511 451
rect 61565 407 61655 451
rect 61709 407 61799 451
rect 61853 407 61943 451
rect 61997 407 62087 451
rect 62141 407 62231 451
rect 62285 407 62500 451
rect -40 343 63 407
rect 62357 343 62500 407
rect -40 299 117 343
rect 171 299 261 343
rect 315 299 405 343
rect 459 299 549 343
rect 603 299 693 343
rect 747 299 837 343
rect 891 299 981 343
rect 1035 299 1125 343
rect 1252 299 1342 343
rect 1396 299 1486 343
rect 1540 299 1630 343
rect 1684 299 1774 343
rect 1828 299 1918 343
rect 1972 299 2062 343
rect 2116 299 2206 343
rect 2260 299 2350 343
rect 2477 299 2567 343
rect 2621 299 2711 343
rect 2765 299 2855 343
rect 2909 299 2999 343
rect 3053 299 3143 343
rect 3197 299 3274 343
rect 60628 299 60718 343
rect 60772 299 60862 343
rect 60916 299 61006 343
rect 61060 299 61150 343
rect 61277 299 61367 343
rect 61421 299 61511 343
rect 61565 299 61655 343
rect 61709 299 61799 343
rect 61853 299 61943 343
rect 61997 299 62087 343
rect 62141 299 62231 343
rect 62285 299 62500 343
rect -40 105 63 299
rect 62357 105 62500 299
rect -40 61 117 105
rect 171 61 261 105
rect 315 61 405 105
rect 459 61 549 105
rect 603 61 693 105
rect 747 61 837 105
rect 891 61 981 105
rect 1035 61 1125 105
rect 1252 61 1342 105
rect 1396 61 1486 105
rect 1540 61 1630 105
rect 1684 61 1774 105
rect 1828 61 1918 105
rect 1972 61 2062 105
rect 2116 61 2206 105
rect 2260 61 2350 105
rect 2477 61 2567 105
rect 2621 61 2711 105
rect 2765 61 2855 105
rect 2909 61 2999 105
rect 3053 61 3143 105
rect 3197 61 3274 105
rect 60628 61 60718 105
rect 60772 61 60862 105
rect 60916 61 61006 105
rect 61060 61 61150 105
rect 61277 61 61367 105
rect 61421 61 61511 105
rect 61565 61 61655 105
rect 61709 61 61799 105
rect 61853 61 61943 105
rect 61997 61 62087 105
rect 62141 61 62231 105
rect 62285 61 62500 105
rect -40 55 63 61
rect 62357 55 62500 61
rect -40 -88 3274 55
rect 60592 -88 62500 55
use sonos_8x8  sonos_8x8_0
array 0 50 1225 0 50 1513
timestamp 1686033482
transform 1 0 0 0 1 0
box -80 -88 1308 1530
<< end >>
