magic
tech sky130A
timestamp 1686033289
<< error_p >>
rect -244 -373 -20 -333
rect -244 -680 96 -373
rect -244 -898 -204 -680
rect -60 -893 96 -680
rect -60 -898 -19 -893
rect -244 -933 -186 -898
rect -222 -943 -186 -933
rect -78 -933 -19 -898
rect -78 -943 -42 -933
rect -222 -961 -204 -943
rect -60 -961 -42 -943
<< dnwell >>
rect -204 -680 -60 -373
rect -204 -893 -59 -680
<< nwell >>
rect -204 -979 -60 -680
<< npd >>
rect -177 -461 -87 -431
<< ndiff >>
rect -177 -389 -87 -381
rect -177 -423 -149 -389
rect -115 -423 -87 -389
rect -177 -431 -87 -423
rect -177 -469 -87 -461
rect -177 -503 -149 -469
rect -115 -503 -87 -469
rect -177 -523 -87 -503
<< ndiffc >>
rect -149 -423 -115 -389
rect -149 -503 -115 -469
<< psubdiff >>
rect -204 -595 -59 -577
rect -204 -629 -149 -595
rect -115 -629 -59 -595
rect -204 -653 -59 -629
<< nsubdiff >>
rect -204 -904 -60 -898
rect -204 -938 -187 -904
rect -77 -938 -60 -904
rect -204 -943 -60 -938
<< psubdiffcont >>
rect -149 -629 -115 -595
<< nsubdiffcont >>
rect -187 -938 -77 -904
<< poly >>
rect -204 -461 -177 -431
rect -87 -461 -60 -431
<< locali >>
rect -154 -389 -44 -373
rect -154 -423 -149 -389
rect -115 -423 -79 -389
rect -45 -423 -44 -389
rect -154 -439 -44 -423
rect -154 -469 -111 -439
rect -154 -503 -149 -469
rect -115 -503 -111 -469
rect -154 -519 -111 -503
rect -204 -629 -149 -595
rect -115 -629 -59 -595
rect -204 -938 -187 -904
rect -77 -938 -60 -904
<< viali >>
rect -79 -423 -45 -389
<< metal1 >>
rect -150 -943 -114 -381
rect -80 -383 -44 -377
rect -85 -389 -39 -383
rect -85 -423 -79 -389
rect -45 -423 -39 -389
rect -85 -429 -39 -423
rect -80 -943 -44 -429
<< end >>
