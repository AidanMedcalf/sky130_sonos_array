magic
tech sky130A
magscale 1 2
timestamp 1685114897
<< error_s >>
rect 492 2709 1094 2747
rect -240 2673 -204 2709
rect -240 2663 -168 2673
rect 492 2663 1128 2709
rect -240 2595 1128 2663
rect -240 2583 -168 2595
rect -240 2573 -204 2583
rect 492 2573 1128 2595
rect -240 2547 1128 2573
rect -204 2358 1094 2547
rect 1152 2494 1346 2530
rect -924 2147 1094 2358
rect 1116 2358 1346 2494
rect 1116 2332 2076 2358
rect -924 1560 1092 2147
rect -1096 1533 1092 1560
rect 1152 1533 2076 2332
rect -1096 1342 0 1533
rect -1060 1306 -898 1342
rect 1152 1335 1992 1533
rect -72 1328 1992 1335
rect -222 1306 1992 1328
rect -1024 1270 -934 1306
rect -1014 970 -946 1270
rect -924 1247 1992 1306
rect -924 1201 1152 1247
rect -924 1172 1180 1201
rect 1224 1190 1235 1230
rect -924 1159 1152 1172
rect -924 1117 1202 1159
rect -924 1102 1224 1117
rect 1456 1102 1648 1104
rect -924 1032 1152 1102
rect 1155 1087 1170 1102
rect -924 972 402 1032
rect 1224 989 1235 1086
rect 1266 1002 1334 1072
rect 1224 988 1256 989
rect 450 972 504 987
rect 594 972 648 987
rect 738 972 792 987
rect 882 972 936 987
rect 1026 972 1080 987
rect -924 970 409 972
rect -1024 965 409 970
rect 450 965 553 972
rect 594 965 697 972
rect 738 965 841 972
rect 882 965 985 972
rect 1026 965 1129 972
rect -1024 948 402 965
rect -1014 942 -946 948
rect -924 942 402 948
rect -1024 920 402 942
rect 466 920 538 957
rect 610 920 682 957
rect 754 920 826 957
rect 898 920 970 957
rect 1042 920 1114 957
rect 1152 923 1202 965
rect 1232 936 1256 988
rect 1266 970 1290 1002
rect 1680 962 1748 994
rect 2098 984 2166 1324
rect 1772 962 2176 984
rect 2098 956 2166 962
rect 1680 924 1748 956
rect 1772 934 2176 956
rect 1152 920 1224 923
rect -1014 834 -946 920
rect -924 910 2076 920
rect 2098 910 2166 934
rect -924 888 2176 910
rect -924 882 2076 888
rect 2098 882 2166 888
rect -924 860 2176 882
rect -924 834 2076 860
rect -1024 812 2076 834
rect -1014 806 -946 812
rect -924 806 2076 812
rect -1024 784 2076 806
rect -1014 760 -946 784
rect -924 774 2076 784
rect 2098 774 2166 860
rect -924 760 2176 774
rect -1024 752 2176 760
rect -1024 746 2076 752
rect 2098 746 2166 752
rect -1024 738 2176 746
rect -1014 732 -946 738
rect -924 732 2176 738
rect -1024 724 2176 732
rect -1024 710 2076 724
rect -1014 624 -946 710
rect -924 638 2076 710
rect 2098 638 2166 724
rect -924 624 2176 638
rect -1024 616 2176 624
rect -1024 610 2076 616
rect 2098 610 2166 616
rect -1024 602 2176 610
rect -1014 596 -946 602
rect -924 596 2176 602
rect -1024 588 2176 596
rect -1024 574 2076 588
rect -1014 488 -946 574
rect -924 564 2076 574
rect 2098 564 2166 588
rect -924 542 2176 564
rect -924 536 2076 542
rect 2098 536 2166 542
rect -924 514 2176 536
rect -924 488 2076 514
rect -1024 466 2076 488
rect -1014 460 -946 466
rect -924 460 2076 466
rect -1024 442 2076 460
rect -1024 438 -620 442
rect -1014 414 -946 438
rect -596 428 -528 442
rect -498 428 2076 442
rect 2098 428 2166 514
rect -1024 392 -620 414
rect -596 392 -528 424
rect -498 406 2176 428
rect -108 400 2076 406
rect 2098 400 2166 406
rect -1014 386 -946 392
rect -1024 364 -620 386
rect -1014 278 -946 364
rect -596 354 -528 386
rect -108 378 2176 400
rect -454 286 -346 288
rect -1024 256 -420 278
rect -182 276 -114 346
rect -108 292 2076 378
rect 2098 292 2166 378
rect -108 270 2176 292
rect -108 264 2076 270
rect 2098 264 2166 270
rect -1014 250 -946 256
rect -1024 228 -420 250
rect -108 242 2176 264
rect -1014 142 -946 228
rect -108 218 2076 242
rect 2098 218 2166 242
rect -108 196 2176 218
rect -108 190 2076 196
rect 2098 190 2166 196
rect -1024 120 -620 142
rect -596 120 -528 152
rect -398 134 -330 170
rect -108 168 2176 190
rect -1014 114 -946 120
rect -1024 92 -620 114
rect -1014 68 -946 92
rect -596 82 -528 114
rect -398 96 -330 132
rect -108 82 2076 168
rect 2098 82 2166 168
rect -1024 46 -620 68
rect -596 46 -528 78
rect -108 60 2176 82
rect -108 54 2076 60
rect 2098 54 2166 60
rect -1014 40 -946 46
rect -1024 18 -620 40
rect -1014 0 -946 18
rect -596 8 -528 40
rect -108 32 2176 54
rect -454 -60 -346 -58
rect -182 -70 -114 0
rect -108 -86 2076 32
rect 2098 0 2166 32
rect -108 -304 2248 -86
rect -108 -312 1224 -304
rect -108 -313 1266 -312
rect -108 -325 1256 -313
rect -108 -333 1224 -325
rect -108 -340 0 -333
rect 2050 -340 2212 -304
rect -138 -519 -114 -497
rect -138 -531 -100 -519
rect -138 -547 -80 -531
rect -150 -552 25 -547
rect -150 -647 -72 -552
rect 10 -562 25 -552
rect -204 -707 -72 -647
rect -150 -724 -72 -707
rect -150 -831 0 -724
rect -124 -876 -100 -831
rect -96 -904 -72 -831
rect -230 -939 0 -930
rect -204 -1090 -203 -939
rect 0 -1090 26 -939
rect -204 -1091 26 -1090
rect 252 -971 1092 -531
rect 252 -1545 1094 -971
rect 1152 -1330 2076 -340
rect 2086 -376 2176 -340
rect 1116 -1356 2076 -1330
rect 1116 -1492 1346 -1356
rect 1152 -1528 1346 -1492
rect -240 -1581 -204 -1545
rect 252 -1571 1128 -1545
rect 1092 -1581 1128 -1571
rect -240 -1593 -168 -1581
rect 1056 -1593 1128 -1581
rect -240 -1661 1128 -1593
rect -240 -1671 -168 -1661
rect 1056 -1671 1128 -1661
rect -240 -1707 -204 -1671
rect 1092 -1707 1128 -1671
<< dnwell >>
rect 0 -32 1 177
<< poly >>
rect 0 100 1 130
rect 0 14 1 58
use sonos_array_corner  sonos_array_corner_0
timestamp 1663090256
transform 1 0 0 0 1 0
box -1096 -1528 276 -156
use sonos_array_corner  sonos_array_corner_1
timestamp 1663090256
transform 1 0 0 0 -1 1002
box -1096 -1528 276 -156
use sonos_array_corner  sonos_array_corner_2
timestamp 1663090256
transform -1 0 1152 0 1 0
box -1096 -1528 276 -156
use sonos_array_corner  sonos_array_corner_3
timestamp 1663090256
transform -1 0 1152 0 -1 1002
box -1096 -1528 276 -156
use sonos_cell  sonos_cell_0
array 0 7 144 0 3 346
timestamp 1684786423
transform 1 0 72 0 1 79
box -224 -332 456 348
use sonos_cell  sonos_cell_1
array 0 7 144 0 3 -346
timestamp 1684786423
transform 1 0 72 0 -1 -115
box -224 -332 456 348
use sonos_endcap_lr  sonos_endcap_lr_0
array 0 0 417 0 3 346
timestamp 1663090256
transform 1 0 0 0 1 0
box -1096 -584 276 776
use sonos_endcap_lr  sonos_endcap_lr_1
array 0 0 417 0 3 346
timestamp 1663090256
transform -1 0 1152 0 -1 1002
box -1096 -584 276 776
use sonos_endcap_tb  sonos_endcap_tb_0
array 0 7 144 0 0 154
timestamp 1663090256
transform 1 0 204 0 1 215
box -568 -1958 792 -586
use sonos_endcap_tb  sonos_endcap_tb_1
array 0 7 144 0 0 -154
timestamp 1663090256
transform 1 0 204 0 -1 787
box -568 -1958 792 -586
<< labels >>
rlabel space -417 -187 -381 -153 1 wl0
rlabel space -417 -113 -381 -79 1 wls0
rlabel space 1533 -93 1569 -59 1 wls0
rlabel space 1533 -161 1569 -127 1 nc0
rlabel space -417 -45 -381 -11 1 nc0
rlabel space -417 23 -381 57 1 wls1
rlabel space 1533 43 1569 77 1 wls1
rlabel space 1533 -25 1569 9 1 nc1
rlabel space -417 91 -381 125 1 nc1
rlabel space 1533 185 1569 219 1 nc2
rlabel space 1533 117 1569 151 1 wl1
rlabel space -417 159 -381 193 1 wl2
rlabel space -417 233 -381 267 1 wls2
rlabel space 1533 253 1569 287 1 wls2
rlabel space 1533 321 1569 355 1 nc3
rlabel space -417 301 -381 335 1 nc2
rlabel space -417 369 -381 403 1 wls3
rlabel space -417 437 -381 471 1 nc3
rlabel space -417 505 -381 539 1 wl4
rlabel space 1533 389 1569 423 1 wls3
rlabel space 1533 463 1569 497 1 wl3
rlabel space 1533 531 1569 565 1 nc4
rlabel space 1533 667 1569 701 1 nc5
rlabel space 1533 877 1569 911 1 nc6
rlabel space 1533 1013 1569 1047 1 nc7
rlabel space 1533 599 1569 633 1 wls4
rlabel space -417 579 -381 613 1 wls4
rlabel space -417 647 -381 681 1 nc4
rlabel space -417 783 -381 817 1 nc5
rlabel space -417 993 -381 1027 1 nc6
rlabel space -417 1129 -381 1163 1 nc7
rlabel space 1533 735 1569 769 1 wls5
rlabel space -417 715 -381 749 1 wls5
rlabel space 1533 809 1569 843 1 wl5
rlabel space -417 851 -381 885 1 wl6
rlabel space 1533 945 1569 979 1 wls6
rlabel space -417 925 -381 959 1 wls6
rlabel space -417 1061 -381 1095 1 wls7
rlabel space 1533 1081 1569 1115 1 wls7
rlabel space 1533 1155 1569 1189 1 wl7
rlabel space 54 -633 90 -597 1 bl0
rlabel space 124 -633 160 -597 1 src0
rlabel space 198 -633 234 -597 1 bl1
rlabel space 268 -633 304 -597 1 src1
rlabel space 342 -633 378 -597 1 bl2
rlabel space 412 -633 448 -597 1 src2
rlabel space 486 -633 522 -597 1 bl3
rlabel space 556 -633 592 -597 1 src3
rlabel space 630 -633 666 -597 1 bl4
rlabel space 700 -633 736 -597 1 src4
rlabel space 774 -633 810 -597 1 bl5
rlabel space 844 -633 880 -597 1 src5
rlabel space 918 -633 954 -597 1 bl6
rlabel space 988 -633 1024 -597 1 src6
rlabel space 1062 -633 1098 -597 1 bl7
rlabel space 1132 -633 1168 -597 1 src7
rlabel space 54 1599 90 1635 1 bl0
rlabel space 124 1599 160 1635 1 src0
rlabel space 198 1599 234 1635 1 bl1
rlabel space 268 1599 304 1635 1 src1
rlabel space 342 1599 378 1635 1 bl2
rlabel space 412 1599 448 1635 1 src2
rlabel space 486 1599 522 1635 1 bl3
rlabel space 556 1599 592 1635 1 src3
rlabel space 630 1599 666 1635 1 bl4
rlabel space 700 1599 736 1635 1 src4
rlabel space 774 1599 810 1635 1 bl5
rlabel space 844 1599 880 1635 1 src5
rlabel space 918 1599 954 1635 1 bl6
rlabel space 988 1599 1024 1635 1 src6
rlabel space 1062 1599 1098 1635 1 bl7
rlabel space 1132 1599 1168 1635 1 src7
rlabel space -111 1382 -50 1440 1 B
rlabel space 1202 1382 1263 1440 1 B
rlabel space 1202 -438 1263 -380 1 B
rlabel space -111 -439 -50 -381 1 B
<< end >>
