magic
tech sky130A
timestamp 1663485803
<< dnwell >>
rect -40 -48 1210 1490
<< psubdiff >>
rect -40 1486 1210 1490
rect -40 1469 0 1486
rect 1173 1469 1210 1486
rect -40 1465 1210 1469
rect -40 1438 -15 1465
rect -40 4 -36 1438
rect -19 4 -15 1438
rect 1185 1438 1210 1465
rect -40 -23 -15 4
rect 1185 4 1189 1438
rect 1206 4 1210 1438
rect 1185 -23 1210 4
rect -40 -27 1210 -23
rect -40 -44 0 -27
rect 1173 -44 1210 -27
rect -40 -48 1210 -44
<< psubdiffcont >>
rect 0 1469 1173 1486
rect -36 4 -19 1438
rect 1189 4 1206 1438
rect 0 -44 1173 -27
<< poly >>
rect 1140 1370 1173 1381
rect 1140 1346 1144 1370
rect 1161 1346 1173 1370
rect 1140 1292 1173 1346
rect 1140 1268 1144 1292
rect 1161 1268 1173 1292
rect 1140 1212 1173 1268
rect 1140 1188 1144 1212
rect 1161 1188 1173 1212
rect 1140 1132 1173 1188
rect 1140 1108 1144 1132
rect 1161 1108 1173 1132
rect 1140 1025 1173 1108
rect 1140 1001 1144 1025
rect 1161 1001 1173 1025
rect 1140 946 1173 1001
rect 1140 922 1144 946
rect 1161 922 1173 946
rect 1140 866 1173 922
rect 1140 842 1144 866
rect 1161 842 1173 866
rect 1140 787 1173 842
rect 1140 763 1144 787
rect 1161 763 1173 787
rect 1140 679 1173 763
rect 1140 655 1144 679
rect 1161 655 1173 679
rect 1140 600 1173 655
rect 1140 576 1144 600
rect 1161 576 1173 600
rect 1140 520 1173 576
rect 1140 496 1144 520
rect 1161 496 1173 520
rect 1140 440 1173 496
rect 1140 416 1144 440
rect 1161 416 1173 440
rect 1140 333 1173 416
rect 1140 309 1144 333
rect 1161 309 1173 333
rect 1140 254 1173 309
rect 1140 230 1144 254
rect 1161 230 1173 254
rect 1140 174 1173 230
rect 1140 150 1144 174
rect 1161 150 1173 174
rect 1140 97 1173 150
rect 1140 73 1144 97
rect 1161 73 1173 97
rect 1140 61 1173 73
<< polycont >>
rect 1144 1346 1161 1370
rect 1144 1268 1161 1292
rect 1144 1188 1161 1212
rect 1144 1108 1161 1132
rect 1144 1001 1161 1025
rect 1144 922 1161 946
rect 1144 842 1161 866
rect 1144 763 1161 787
rect 1144 655 1161 679
rect 1144 576 1161 600
rect 1144 496 1161 520
rect 1144 416 1161 440
rect 1144 309 1161 333
rect 1144 230 1161 254
rect 1144 150 1161 174
rect 1144 73 1161 97
<< locali >>
rect -36 1469 0 1486
rect 1173 1469 1206 1486
rect -36 1438 -19 1469
rect 39 1438 1113 1469
rect 1189 1438 1206 1469
rect 1136 1370 1189 1381
rect 1136 1346 1144 1370
rect 1161 1346 1189 1370
rect -19 1312 0 1346
rect 1136 1292 1189 1346
rect 1136 1268 1144 1292
rect 1161 1268 1189 1292
rect 1136 1212 1189 1268
rect 1136 1188 1144 1212
rect 1161 1188 1189 1212
rect -19 1134 0 1168
rect 1136 1132 1189 1188
rect 1136 1108 1144 1132
rect 1161 1108 1189 1132
rect 1136 1025 1189 1108
rect 1136 1001 1144 1025
rect 1161 1001 1189 1025
rect -19 966 0 1000
rect 1136 946 1189 1001
rect 1136 922 1144 946
rect 1161 922 1189 946
rect 1136 866 1189 922
rect 1136 842 1144 866
rect 1161 842 1189 866
rect -19 788 0 822
rect 1136 787 1189 842
rect 1136 763 1144 787
rect 1161 763 1189 787
rect 1136 679 1189 763
rect 1136 655 1144 679
rect 1161 655 1189 679
rect -19 620 0 654
rect 1136 600 1189 655
rect 1136 576 1144 600
rect 1161 576 1189 600
rect 1136 520 1189 576
rect 1136 496 1144 520
rect 1161 496 1189 520
rect -19 442 0 476
rect 1136 440 1189 496
rect 1136 416 1144 440
rect 1161 416 1189 440
rect 1136 333 1189 416
rect 1136 309 1144 333
rect 1161 309 1189 333
rect -19 274 0 308
rect 1136 254 1189 309
rect 1136 230 1144 254
rect 1161 230 1189 254
rect 1136 174 1189 230
rect 1136 150 1144 174
rect 1161 150 1189 174
rect -19 96 0 130
rect 1136 97 1189 150
rect 1136 73 1144 97
rect 1161 73 1189 97
rect 1136 61 1189 73
rect -36 -27 -19 4
rect 39 -27 1113 4
rect 1189 -27 1206 4
rect -36 -44 0 -27
rect 1173 -44 1206 -27
<< metal1 >>
rect 95 1390 1152 1436
rect 92 6 1155 52
use sonos_cell_mirrored  sonos_cell_mirrored_0
array 0 7 144 0 3 346
timestamp 1663485803
transform 1 0 -80 0 1 -80
box 80 80 380 484
<< end >>
