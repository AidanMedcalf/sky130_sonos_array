magic
tech sky130A
magscale 1 2
timestamp 1684788722
<< error_s >>
rect 243214 296750 243394 296838
rect 243502 296750 243682 296838
rect 243790 296750 243970 296838
rect 244078 296750 244258 296838
rect 244366 296750 244546 296838
rect 244654 296750 244834 296838
rect 244942 296750 245122 296838
rect 245230 296750 245410 296838
rect 245664 296750 245844 296838
rect 245952 296750 246132 296838
rect 246240 296750 246420 296838
rect 246528 296750 246708 296838
rect 246816 296750 246996 296838
rect 247104 296750 247284 296838
rect 247392 296750 247572 296838
rect 247680 296750 247860 296838
rect 248114 296750 248294 296838
rect 248402 296750 248582 296838
rect 248690 296750 248870 296838
rect 248978 296750 249158 296838
rect 249266 296750 249446 296838
rect 249554 296750 249734 296838
rect 249842 296750 250022 296838
rect 250130 296750 250310 296838
rect 250564 296750 250744 296838
rect 250852 296750 251032 296838
rect 251140 296750 251320 296838
rect 251428 296750 251608 296838
rect 251716 296750 251896 296838
rect 252004 296750 252184 296838
rect 252292 296750 252472 296838
rect 252580 296750 252760 296838
rect 253014 296750 253194 296838
rect 253302 296750 253482 296838
rect 253590 296750 253770 296838
rect 253878 296750 254058 296838
rect 254166 296750 254346 296838
rect 254454 296750 254634 296838
rect 254742 296750 254922 296838
rect 255030 296750 255210 296838
rect 255464 296750 255644 296838
rect 255752 296750 255932 296838
rect 256040 296750 256220 296838
rect 256328 296750 256508 296838
rect 256616 296750 256796 296838
rect 256904 296750 257084 296838
rect 257192 296750 257372 296838
rect 257480 296750 257660 296838
rect 257914 296750 258094 296838
rect 258202 296750 258382 296838
rect 258490 296750 258670 296838
rect 258778 296750 258958 296838
rect 259066 296750 259246 296838
rect 259354 296750 259534 296838
rect 259642 296750 259822 296838
rect 259930 296750 260110 296838
rect 260364 296750 260544 296838
rect 260652 296750 260832 296838
rect 260940 296750 261120 296838
rect 261228 296750 261408 296838
rect 261516 296750 261696 296838
rect 261804 296750 261984 296838
rect 262092 296750 262272 296838
rect 262380 296750 262560 296838
rect 262814 296750 262994 296838
rect 263102 296750 263282 296838
rect 263390 296750 263570 296838
rect 263678 296750 263858 296838
rect 263966 296750 264146 296838
rect 264254 296750 264434 296838
rect 264542 296750 264722 296838
rect 264830 296750 265010 296838
rect 265264 296750 265444 296838
rect 265552 296750 265732 296838
rect 265840 296750 266020 296838
rect 266128 296750 266308 296838
rect 266416 296750 266596 296838
rect 266704 296750 266884 296838
rect 266992 296750 267172 296838
rect 267280 296750 267460 296838
rect 267714 296750 267894 296838
rect 268002 296750 268182 296838
rect 268290 296750 268470 296838
rect 268578 296750 268758 296838
rect 268866 296750 269046 296838
rect 269154 296750 269334 296838
rect 269442 296750 269622 296838
rect 269730 296750 269910 296838
rect 270164 296750 270344 296838
rect 270452 296750 270632 296838
rect 270740 296750 270920 296838
rect 271028 296750 271208 296838
rect 271316 296750 271496 296838
rect 271604 296750 271784 296838
rect 271892 296750 272072 296838
rect 272180 296750 272360 296838
rect 272614 296750 272794 296838
rect 272902 296750 273082 296838
rect 273190 296750 273370 296838
rect 273478 296750 273658 296838
rect 273766 296750 273946 296838
rect 274054 296750 274234 296838
rect 274342 296750 274522 296838
rect 274630 296750 274810 296838
rect 275064 296750 275244 296838
rect 275352 296750 275532 296838
rect 275640 296750 275820 296838
rect 275928 296750 276108 296838
rect 276216 296750 276396 296838
rect 276504 296750 276684 296838
rect 276792 296750 276972 296838
rect 277080 296750 277260 296838
rect 277514 296750 277694 296838
rect 277802 296750 277982 296838
rect 278090 296750 278270 296838
rect 278378 296750 278558 296838
rect 278666 296750 278846 296838
rect 278954 296750 279134 296838
rect 279242 296750 279422 296838
rect 279530 296750 279710 296838
rect 279964 296750 280144 296838
rect 280252 296750 280432 296838
rect 280540 296750 280720 296838
rect 280828 296750 281008 296838
rect 281116 296750 281296 296838
rect 281404 296750 281584 296838
rect 281692 296750 281872 296838
rect 281980 296750 282160 296838
rect 282414 296750 282594 296838
rect 282702 296750 282882 296838
rect 282990 296750 283170 296838
rect 283278 296750 283458 296838
rect 283566 296750 283746 296838
rect 283854 296750 284034 296838
rect 284142 296750 284322 296838
rect 284430 296750 284610 296838
rect 284864 296750 285044 296838
rect 285152 296750 285332 296838
rect 285440 296750 285620 296838
rect 285728 296750 285908 296838
rect 286016 296750 286196 296838
rect 286304 296750 286484 296838
rect 286592 296750 286772 296838
rect 286880 296750 287060 296838
rect 287314 296750 287494 296838
rect 287602 296750 287782 296838
rect 287890 296750 288070 296838
rect 288178 296750 288358 296838
rect 288466 296750 288646 296838
rect 288754 296750 288934 296838
rect 289042 296750 289222 296838
rect 289330 296750 289510 296838
rect 289764 296750 289944 296838
rect 290052 296750 290232 296838
rect 290340 296750 290520 296838
rect 290628 296750 290808 296838
rect 290916 296750 291096 296838
rect 291204 296750 291384 296838
rect 291492 296750 291672 296838
rect 291780 296750 291960 296838
rect 292214 296750 292394 296838
rect 292502 296750 292682 296838
rect 292790 296750 292970 296838
rect 293078 296750 293258 296838
rect 293366 296750 293546 296838
rect 293654 296750 293834 296838
rect 293942 296750 294122 296838
rect 294230 296750 294410 296838
rect 294664 296750 294844 296838
rect 294952 296750 295132 296838
rect 295240 296750 295420 296838
rect 295528 296750 295708 296838
rect 295816 296750 295996 296838
rect 296104 296750 296284 296838
rect 296392 296750 296572 296838
rect 296680 296750 296860 296838
rect 297114 296750 297294 296838
rect 297402 296750 297582 296838
rect 297690 296750 297870 296838
rect 297978 296750 298158 296838
rect 298266 296750 298446 296838
rect 298554 296750 298734 296838
rect 298842 296750 299022 296838
rect 299130 296750 299310 296838
rect 299564 296750 299744 296838
rect 299852 296750 300032 296838
rect 300140 296750 300320 296838
rect 300428 296750 300608 296838
rect 300716 296750 300896 296838
rect 301004 296750 301184 296838
rect 301292 296750 301472 296838
rect 301580 296750 301760 296838
rect 302014 296750 302194 296838
rect 302302 296750 302482 296838
rect 302590 296750 302770 296838
rect 302878 296750 303058 296838
rect 303166 296750 303346 296838
rect 303454 296750 303634 296838
rect 303742 296750 303922 296838
rect 304030 296750 304210 296838
rect 304464 296750 304644 296838
rect 304752 296750 304932 296838
rect 305040 296750 305220 296838
rect 305328 296750 305508 296838
rect 305616 296750 305796 296838
rect 305904 296750 306084 296838
rect 306192 296750 306372 296838
rect 306480 296750 306660 296838
rect 306914 296750 307094 296838
rect 307202 296750 307382 296838
rect 307490 296750 307670 296838
rect 307778 296750 307958 296838
rect 308066 296750 308246 296838
rect 308354 296750 308534 296838
rect 308642 296750 308822 296838
rect 308930 296750 309110 296838
rect 309364 296750 309544 296838
rect 309652 296750 309832 296838
rect 309940 296750 310120 296838
rect 310228 296750 310408 296838
rect 310516 296750 310696 296838
rect 310804 296750 310984 296838
rect 311092 296750 311272 296838
rect 311380 296750 311560 296838
rect 311814 296750 311994 296838
rect 312102 296750 312282 296838
rect 312390 296750 312570 296838
rect 312678 296750 312858 296838
rect 312966 296750 313146 296838
rect 313254 296750 313434 296838
rect 313542 296750 313722 296838
rect 313830 296750 314010 296838
rect 314264 296750 314444 296838
rect 314552 296750 314732 296838
rect 314840 296750 315020 296838
rect 315128 296750 315308 296838
rect 315416 296750 315596 296838
rect 315704 296750 315884 296838
rect 315992 296750 316172 296838
rect 316280 296750 316460 296838
rect 316714 296750 316894 296838
rect 317002 296750 317182 296838
rect 317290 296750 317470 296838
rect 317578 296750 317758 296838
rect 317866 296750 318046 296838
rect 318154 296750 318334 296838
rect 318442 296750 318622 296838
rect 318730 296750 318910 296838
rect 319164 296750 319344 296838
rect 319452 296750 319632 296838
rect 319740 296750 319920 296838
rect 320028 296750 320208 296838
rect 320316 296750 320496 296838
rect 320604 296750 320784 296838
rect 320892 296750 321072 296838
rect 321180 296750 321360 296838
rect 321614 296750 321794 296838
rect 321902 296750 322082 296838
rect 322190 296750 322370 296838
rect 322478 296750 322658 296838
rect 322766 296750 322946 296838
rect 323054 296750 323234 296838
rect 323342 296750 323522 296838
rect 323630 296750 323810 296838
rect 324064 296750 324244 296838
rect 324352 296750 324532 296838
rect 324640 296750 324820 296838
rect 324928 296750 325108 296838
rect 325216 296750 325396 296838
rect 325504 296750 325684 296838
rect 325792 296750 325972 296838
rect 326080 296750 326260 296838
rect 326514 296750 326694 296838
rect 326802 296750 326982 296838
rect 327090 296750 327270 296838
rect 327378 296750 327558 296838
rect 327666 296750 327846 296838
rect 327954 296750 328134 296838
rect 328242 296750 328422 296838
rect 328530 296750 328710 296838
rect 328964 296750 329144 296838
rect 329252 296750 329432 296838
rect 329540 296750 329720 296838
rect 329828 296750 330008 296838
rect 330116 296750 330296 296838
rect 330404 296750 330584 296838
rect 330692 296750 330872 296838
rect 330980 296750 331160 296838
rect 331414 296750 331594 296838
rect 331702 296750 331882 296838
rect 331990 296750 332170 296838
rect 332278 296750 332458 296838
rect 332566 296750 332746 296838
rect 332854 296750 333034 296838
rect 333142 296750 333322 296838
rect 333430 296750 333610 296838
rect 333864 296750 334044 296838
rect 334152 296750 334332 296838
rect 334440 296750 334620 296838
rect 334728 296750 334908 296838
rect 335016 296750 335196 296838
rect 335304 296750 335484 296838
rect 335592 296750 335772 296838
rect 335880 296750 336060 296838
rect 336314 296750 336494 296838
rect 336602 296750 336782 296838
rect 336890 296750 337070 296838
rect 337178 296750 337358 296838
rect 337466 296750 337646 296838
rect 337754 296750 337934 296838
rect 338042 296750 338222 296838
rect 338330 296750 338510 296838
rect 338764 296750 338944 296838
rect 339052 296750 339232 296838
rect 339340 296750 339520 296838
rect 339628 296750 339808 296838
rect 339916 296750 340096 296838
rect 340204 296750 340384 296838
rect 340492 296750 340672 296838
rect 340780 296750 340960 296838
rect 341214 296750 341394 296838
rect 341502 296750 341682 296838
rect 341790 296750 341970 296838
rect 342078 296750 342258 296838
rect 342366 296750 342546 296838
rect 342654 296750 342834 296838
rect 342942 296750 343122 296838
rect 343230 296750 343410 296838
rect 343664 296750 343844 296838
rect 343952 296750 344132 296838
rect 344240 296750 344420 296838
rect 344528 296750 344708 296838
rect 344816 296750 344996 296838
rect 345104 296750 345284 296838
rect 345392 296750 345572 296838
rect 345680 296750 345860 296838
rect 346114 296750 346294 296838
rect 346402 296750 346582 296838
rect 346690 296750 346870 296838
rect 346978 296750 347158 296838
rect 347266 296750 347446 296838
rect 347554 296750 347734 296838
rect 347842 296750 348022 296838
rect 348130 296750 348310 296838
rect 348564 296750 348744 296838
rect 348852 296750 349032 296838
rect 349140 296750 349320 296838
rect 349428 296750 349608 296838
rect 349716 296750 349896 296838
rect 350004 296750 350184 296838
rect 350292 296750 350472 296838
rect 350580 296750 350760 296838
rect 351014 296750 351194 296838
rect 351302 296750 351482 296838
rect 351590 296750 351770 296838
rect 351878 296750 352058 296838
rect 352166 296750 352346 296838
rect 352454 296750 352634 296838
rect 352742 296750 352922 296838
rect 353030 296750 353210 296838
rect 353464 296750 353644 296838
rect 353752 296750 353932 296838
rect 354040 296750 354220 296838
rect 354328 296750 354508 296838
rect 354616 296750 354796 296838
rect 354904 296750 355084 296838
rect 355192 296750 355372 296838
rect 355480 296750 355660 296838
rect 355914 296750 356094 296838
rect 356202 296750 356382 296838
rect 356490 296750 356670 296838
rect 356778 296750 356958 296838
rect 357066 296750 357246 296838
rect 357354 296750 357534 296838
rect 357642 296750 357822 296838
rect 357930 296750 358110 296838
rect 358364 296750 358544 296838
rect 358652 296750 358832 296838
rect 358940 296750 359120 296838
rect 359228 296750 359408 296838
rect 359516 296750 359696 296838
rect 359804 296750 359984 296838
rect 360092 296750 360272 296838
rect 360380 296750 360560 296838
rect 360814 296750 360994 296838
rect 361102 296750 361282 296838
rect 361390 296750 361570 296838
rect 361678 296750 361858 296838
rect 361966 296750 362146 296838
rect 362254 296750 362434 296838
rect 362542 296750 362722 296838
rect 362830 296750 363010 296838
rect 363264 296750 363444 296838
rect 363552 296750 363732 296838
rect 363840 296750 364020 296838
rect 364128 296750 364308 296838
rect 364416 296750 364596 296838
rect 364704 296750 364884 296838
rect 364992 296750 365172 296838
rect 365280 296750 365460 296838
rect 365714 296750 365894 296838
rect 366002 296750 366182 296838
rect 366290 296750 366470 296838
rect 366578 296750 366758 296838
rect 366866 296750 367046 296838
rect 367154 296750 367334 296838
rect 367442 296750 367622 296838
rect 367730 296750 367910 296838
rect 243214 296274 243394 296362
rect 243502 296274 243682 296362
rect 243790 296274 243970 296362
rect 244078 296274 244258 296362
rect 244366 296274 244546 296362
rect 244654 296274 244834 296362
rect 244942 296274 245122 296362
rect 245230 296274 245410 296362
rect 245664 296274 245844 296362
rect 245952 296274 246132 296362
rect 246240 296274 246420 296362
rect 246528 296274 246708 296362
rect 246816 296274 246996 296362
rect 247104 296274 247284 296362
rect 247392 296274 247572 296362
rect 247680 296274 247860 296362
rect 248114 296274 248294 296362
rect 248402 296274 248582 296362
rect 248690 296274 248870 296362
rect 248978 296274 249158 296362
rect 249266 296274 249446 296362
rect 249554 296274 249734 296362
rect 249842 296274 250022 296362
rect 250130 296274 250310 296362
rect 250564 296274 250744 296362
rect 250852 296274 251032 296362
rect 251140 296274 251320 296362
rect 251428 296274 251608 296362
rect 251716 296274 251896 296362
rect 252004 296274 252184 296362
rect 252292 296274 252472 296362
rect 252580 296274 252760 296362
rect 253014 296274 253194 296362
rect 253302 296274 253482 296362
rect 253590 296274 253770 296362
rect 253878 296274 254058 296362
rect 254166 296274 254346 296362
rect 254454 296274 254634 296362
rect 254742 296274 254922 296362
rect 255030 296274 255210 296362
rect 255464 296274 255644 296362
rect 255752 296274 255932 296362
rect 256040 296274 256220 296362
rect 256328 296274 256508 296362
rect 256616 296274 256796 296362
rect 256904 296274 257084 296362
rect 257192 296274 257372 296362
rect 257480 296274 257660 296362
rect 257914 296274 258094 296362
rect 258202 296274 258382 296362
rect 258490 296274 258670 296362
rect 258778 296274 258958 296362
rect 259066 296274 259246 296362
rect 259354 296274 259534 296362
rect 259642 296274 259822 296362
rect 259930 296274 260110 296362
rect 260364 296274 260544 296362
rect 260652 296274 260832 296362
rect 260940 296274 261120 296362
rect 261228 296274 261408 296362
rect 261516 296274 261696 296362
rect 261804 296274 261984 296362
rect 262092 296274 262272 296362
rect 262380 296274 262560 296362
rect 262814 296274 262994 296362
rect 263102 296274 263282 296362
rect 263390 296274 263570 296362
rect 263678 296274 263858 296362
rect 263966 296274 264146 296362
rect 264254 296274 264434 296362
rect 264542 296274 264722 296362
rect 264830 296274 265010 296362
rect 265264 296274 265444 296362
rect 265552 296274 265732 296362
rect 265840 296274 266020 296362
rect 266128 296274 266308 296362
rect 266416 296274 266596 296362
rect 266704 296274 266884 296362
rect 266992 296274 267172 296362
rect 267280 296274 267460 296362
rect 267714 296274 267894 296362
rect 268002 296274 268182 296362
rect 268290 296274 268470 296362
rect 268578 296274 268758 296362
rect 268866 296274 269046 296362
rect 269154 296274 269334 296362
rect 269442 296274 269622 296362
rect 269730 296274 269910 296362
rect 270164 296274 270344 296362
rect 270452 296274 270632 296362
rect 270740 296274 270920 296362
rect 271028 296274 271208 296362
rect 271316 296274 271496 296362
rect 271604 296274 271784 296362
rect 271892 296274 272072 296362
rect 272180 296274 272360 296362
rect 272614 296274 272794 296362
rect 272902 296274 273082 296362
rect 273190 296274 273370 296362
rect 273478 296274 273658 296362
rect 273766 296274 273946 296362
rect 274054 296274 274234 296362
rect 274342 296274 274522 296362
rect 274630 296274 274810 296362
rect 275064 296274 275244 296362
rect 275352 296274 275532 296362
rect 275640 296274 275820 296362
rect 275928 296274 276108 296362
rect 276216 296274 276396 296362
rect 276504 296274 276684 296362
rect 276792 296274 276972 296362
rect 277080 296274 277260 296362
rect 277514 296274 277694 296362
rect 277802 296274 277982 296362
rect 278090 296274 278270 296362
rect 278378 296274 278558 296362
rect 278666 296274 278846 296362
rect 278954 296274 279134 296362
rect 279242 296274 279422 296362
rect 279530 296274 279710 296362
rect 279964 296274 280144 296362
rect 280252 296274 280432 296362
rect 280540 296274 280720 296362
rect 280828 296274 281008 296362
rect 281116 296274 281296 296362
rect 281404 296274 281584 296362
rect 281692 296274 281872 296362
rect 281980 296274 282160 296362
rect 282414 296274 282594 296362
rect 282702 296274 282882 296362
rect 282990 296274 283170 296362
rect 283278 296274 283458 296362
rect 283566 296274 283746 296362
rect 283854 296274 284034 296362
rect 284142 296274 284322 296362
rect 284430 296274 284610 296362
rect 284864 296274 285044 296362
rect 285152 296274 285332 296362
rect 285440 296274 285620 296362
rect 285728 296274 285908 296362
rect 286016 296274 286196 296362
rect 286304 296274 286484 296362
rect 286592 296274 286772 296362
rect 286880 296274 287060 296362
rect 287314 296274 287494 296362
rect 287602 296274 287782 296362
rect 287890 296274 288070 296362
rect 288178 296274 288358 296362
rect 288466 296274 288646 296362
rect 288754 296274 288934 296362
rect 289042 296274 289222 296362
rect 289330 296274 289510 296362
rect 289764 296274 289944 296362
rect 290052 296274 290232 296362
rect 290340 296274 290520 296362
rect 290628 296274 290808 296362
rect 290916 296274 291096 296362
rect 291204 296274 291384 296362
rect 291492 296274 291672 296362
rect 291780 296274 291960 296362
rect 292214 296274 292394 296362
rect 292502 296274 292682 296362
rect 292790 296274 292970 296362
rect 293078 296274 293258 296362
rect 293366 296274 293546 296362
rect 293654 296274 293834 296362
rect 293942 296274 294122 296362
rect 294230 296274 294410 296362
rect 294664 296274 294844 296362
rect 294952 296274 295132 296362
rect 295240 296274 295420 296362
rect 295528 296274 295708 296362
rect 295816 296274 295996 296362
rect 296104 296274 296284 296362
rect 296392 296274 296572 296362
rect 296680 296274 296860 296362
rect 297114 296274 297294 296362
rect 297402 296274 297582 296362
rect 297690 296274 297870 296362
rect 297978 296274 298158 296362
rect 298266 296274 298446 296362
rect 298554 296274 298734 296362
rect 298842 296274 299022 296362
rect 299130 296274 299310 296362
rect 299564 296274 299744 296362
rect 299852 296274 300032 296362
rect 300140 296274 300320 296362
rect 300428 296274 300608 296362
rect 300716 296274 300896 296362
rect 301004 296274 301184 296362
rect 301292 296274 301472 296362
rect 301580 296274 301760 296362
rect 302014 296274 302194 296362
rect 302302 296274 302482 296362
rect 302590 296274 302770 296362
rect 302878 296274 303058 296362
rect 303166 296274 303346 296362
rect 303454 296274 303634 296362
rect 303742 296274 303922 296362
rect 304030 296274 304210 296362
rect 304464 296274 304644 296362
rect 304752 296274 304932 296362
rect 305040 296274 305220 296362
rect 305328 296274 305508 296362
rect 305616 296274 305796 296362
rect 305904 296274 306084 296362
rect 306192 296274 306372 296362
rect 306480 296274 306660 296362
rect 306914 296274 307094 296362
rect 307202 296274 307382 296362
rect 307490 296274 307670 296362
rect 307778 296274 307958 296362
rect 308066 296274 308246 296362
rect 308354 296274 308534 296362
rect 308642 296274 308822 296362
rect 308930 296274 309110 296362
rect 309364 296274 309544 296362
rect 309652 296274 309832 296362
rect 309940 296274 310120 296362
rect 310228 296274 310408 296362
rect 310516 296274 310696 296362
rect 310804 296274 310984 296362
rect 311092 296274 311272 296362
rect 311380 296274 311560 296362
rect 311814 296274 311994 296362
rect 312102 296274 312282 296362
rect 312390 296274 312570 296362
rect 312678 296274 312858 296362
rect 312966 296274 313146 296362
rect 313254 296274 313434 296362
rect 313542 296274 313722 296362
rect 313830 296274 314010 296362
rect 314264 296274 314444 296362
rect 314552 296274 314732 296362
rect 314840 296274 315020 296362
rect 315128 296274 315308 296362
rect 315416 296274 315596 296362
rect 315704 296274 315884 296362
rect 315992 296274 316172 296362
rect 316280 296274 316460 296362
rect 316714 296274 316894 296362
rect 317002 296274 317182 296362
rect 317290 296274 317470 296362
rect 317578 296274 317758 296362
rect 317866 296274 318046 296362
rect 318154 296274 318334 296362
rect 318442 296274 318622 296362
rect 318730 296274 318910 296362
rect 319164 296274 319344 296362
rect 319452 296274 319632 296362
rect 319740 296274 319920 296362
rect 320028 296274 320208 296362
rect 320316 296274 320496 296362
rect 320604 296274 320784 296362
rect 320892 296274 321072 296362
rect 321180 296274 321360 296362
rect 321614 296274 321794 296362
rect 321902 296274 322082 296362
rect 322190 296274 322370 296362
rect 322478 296274 322658 296362
rect 322766 296274 322946 296362
rect 323054 296274 323234 296362
rect 323342 296274 323522 296362
rect 323630 296274 323810 296362
rect 324064 296274 324244 296362
rect 324352 296274 324532 296362
rect 324640 296274 324820 296362
rect 324928 296274 325108 296362
rect 325216 296274 325396 296362
rect 325504 296274 325684 296362
rect 325792 296274 325972 296362
rect 326080 296274 326260 296362
rect 326514 296274 326694 296362
rect 326802 296274 326982 296362
rect 327090 296274 327270 296362
rect 327378 296274 327558 296362
rect 327666 296274 327846 296362
rect 327954 296274 328134 296362
rect 328242 296274 328422 296362
rect 328530 296274 328710 296362
rect 328964 296274 329144 296362
rect 329252 296274 329432 296362
rect 329540 296274 329720 296362
rect 329828 296274 330008 296362
rect 330116 296274 330296 296362
rect 330404 296274 330584 296362
rect 330692 296274 330872 296362
rect 330980 296274 331160 296362
rect 331414 296274 331594 296362
rect 331702 296274 331882 296362
rect 331990 296274 332170 296362
rect 332278 296274 332458 296362
rect 332566 296274 332746 296362
rect 332854 296274 333034 296362
rect 333142 296274 333322 296362
rect 333430 296274 333610 296362
rect 333864 296274 334044 296362
rect 334152 296274 334332 296362
rect 334440 296274 334620 296362
rect 334728 296274 334908 296362
rect 335016 296274 335196 296362
rect 335304 296274 335484 296362
rect 335592 296274 335772 296362
rect 335880 296274 336060 296362
rect 336314 296274 336494 296362
rect 336602 296274 336782 296362
rect 336890 296274 337070 296362
rect 337178 296274 337358 296362
rect 337466 296274 337646 296362
rect 337754 296274 337934 296362
rect 338042 296274 338222 296362
rect 338330 296274 338510 296362
rect 338764 296274 338944 296362
rect 339052 296274 339232 296362
rect 339340 296274 339520 296362
rect 339628 296274 339808 296362
rect 339916 296274 340096 296362
rect 340204 296274 340384 296362
rect 340492 296274 340672 296362
rect 340780 296274 340960 296362
rect 341214 296274 341394 296362
rect 341502 296274 341682 296362
rect 341790 296274 341970 296362
rect 342078 296274 342258 296362
rect 342366 296274 342546 296362
rect 342654 296274 342834 296362
rect 342942 296274 343122 296362
rect 343230 296274 343410 296362
rect 343664 296274 343844 296362
rect 343952 296274 344132 296362
rect 344240 296274 344420 296362
rect 344528 296274 344708 296362
rect 344816 296274 344996 296362
rect 345104 296274 345284 296362
rect 345392 296274 345572 296362
rect 345680 296274 345860 296362
rect 346114 296274 346294 296362
rect 346402 296274 346582 296362
rect 346690 296274 346870 296362
rect 346978 296274 347158 296362
rect 347266 296274 347446 296362
rect 347554 296274 347734 296362
rect 347842 296274 348022 296362
rect 348130 296274 348310 296362
rect 348564 296274 348744 296362
rect 348852 296274 349032 296362
rect 349140 296274 349320 296362
rect 349428 296274 349608 296362
rect 349716 296274 349896 296362
rect 350004 296274 350184 296362
rect 350292 296274 350472 296362
rect 350580 296274 350760 296362
rect 351014 296274 351194 296362
rect 351302 296274 351482 296362
rect 351590 296274 351770 296362
rect 351878 296274 352058 296362
rect 352166 296274 352346 296362
rect 352454 296274 352634 296362
rect 352742 296274 352922 296362
rect 353030 296274 353210 296362
rect 353464 296274 353644 296362
rect 353752 296274 353932 296362
rect 354040 296274 354220 296362
rect 354328 296274 354508 296362
rect 354616 296274 354796 296362
rect 354904 296274 355084 296362
rect 355192 296274 355372 296362
rect 355480 296274 355660 296362
rect 355914 296274 356094 296362
rect 356202 296274 356382 296362
rect 356490 296274 356670 296362
rect 356778 296274 356958 296362
rect 357066 296274 357246 296362
rect 357354 296274 357534 296362
rect 357642 296274 357822 296362
rect 357930 296274 358110 296362
rect 358364 296274 358544 296362
rect 358652 296274 358832 296362
rect 358940 296274 359120 296362
rect 359228 296274 359408 296362
rect 359516 296274 359696 296362
rect 359804 296274 359984 296362
rect 360092 296274 360272 296362
rect 360380 296274 360560 296362
rect 360814 296274 360994 296362
rect 361102 296274 361282 296362
rect 361390 296274 361570 296362
rect 361678 296274 361858 296362
rect 361966 296274 362146 296362
rect 362254 296274 362434 296362
rect 362542 296274 362722 296362
rect 362830 296274 363010 296362
rect 363264 296274 363444 296362
rect 363552 296274 363732 296362
rect 363840 296274 364020 296362
rect 364128 296274 364308 296362
rect 364416 296274 364596 296362
rect 364704 296274 364884 296362
rect 364992 296274 365172 296362
rect 365280 296274 365460 296362
rect 365714 296274 365894 296362
rect 366002 296274 366182 296362
rect 366290 296274 366470 296362
rect 366578 296274 366758 296362
rect 366866 296274 367046 296362
rect 367154 296274 367334 296362
rect 367442 296274 367622 296362
rect 367730 296274 367910 296362
rect 243214 296058 243394 296146
rect 243502 296058 243682 296146
rect 243790 296058 243970 296146
rect 244078 296058 244258 296146
rect 244366 296058 244546 296146
rect 244654 296058 244834 296146
rect 244942 296058 245122 296146
rect 245230 296058 245410 296146
rect 245664 296058 245844 296146
rect 245952 296058 246132 296146
rect 246240 296058 246420 296146
rect 246528 296058 246708 296146
rect 246816 296058 246996 296146
rect 247104 296058 247284 296146
rect 247392 296058 247572 296146
rect 247680 296058 247860 296146
rect 248114 296058 248294 296146
rect 248402 296058 248582 296146
rect 248690 296058 248870 296146
rect 248978 296058 249158 296146
rect 249266 296058 249446 296146
rect 249554 296058 249734 296146
rect 249842 296058 250022 296146
rect 250130 296058 250310 296146
rect 250564 296058 250744 296146
rect 250852 296058 251032 296146
rect 251140 296058 251320 296146
rect 251428 296058 251608 296146
rect 251716 296058 251896 296146
rect 252004 296058 252184 296146
rect 252292 296058 252472 296146
rect 252580 296058 252760 296146
rect 253014 296058 253194 296146
rect 253302 296058 253482 296146
rect 253590 296058 253770 296146
rect 253878 296058 254058 296146
rect 254166 296058 254346 296146
rect 254454 296058 254634 296146
rect 254742 296058 254922 296146
rect 255030 296058 255210 296146
rect 255464 296058 255644 296146
rect 255752 296058 255932 296146
rect 256040 296058 256220 296146
rect 256328 296058 256508 296146
rect 256616 296058 256796 296146
rect 256904 296058 257084 296146
rect 257192 296058 257372 296146
rect 257480 296058 257660 296146
rect 257914 296058 258094 296146
rect 258202 296058 258382 296146
rect 258490 296058 258670 296146
rect 258778 296058 258958 296146
rect 259066 296058 259246 296146
rect 259354 296058 259534 296146
rect 259642 296058 259822 296146
rect 259930 296058 260110 296146
rect 260364 296058 260544 296146
rect 260652 296058 260832 296146
rect 260940 296058 261120 296146
rect 261228 296058 261408 296146
rect 261516 296058 261696 296146
rect 261804 296058 261984 296146
rect 262092 296058 262272 296146
rect 262380 296058 262560 296146
rect 262814 296058 262994 296146
rect 263102 296058 263282 296146
rect 263390 296058 263570 296146
rect 263678 296058 263858 296146
rect 263966 296058 264146 296146
rect 264254 296058 264434 296146
rect 264542 296058 264722 296146
rect 264830 296058 265010 296146
rect 265264 296058 265444 296146
rect 265552 296058 265732 296146
rect 265840 296058 266020 296146
rect 266128 296058 266308 296146
rect 266416 296058 266596 296146
rect 266704 296058 266884 296146
rect 266992 296058 267172 296146
rect 267280 296058 267460 296146
rect 267714 296058 267894 296146
rect 268002 296058 268182 296146
rect 268290 296058 268470 296146
rect 268578 296058 268758 296146
rect 268866 296058 269046 296146
rect 269154 296058 269334 296146
rect 269442 296058 269622 296146
rect 269730 296058 269910 296146
rect 270164 296058 270344 296146
rect 270452 296058 270632 296146
rect 270740 296058 270920 296146
rect 271028 296058 271208 296146
rect 271316 296058 271496 296146
rect 271604 296058 271784 296146
rect 271892 296058 272072 296146
rect 272180 296058 272360 296146
rect 272614 296058 272794 296146
rect 272902 296058 273082 296146
rect 273190 296058 273370 296146
rect 273478 296058 273658 296146
rect 273766 296058 273946 296146
rect 274054 296058 274234 296146
rect 274342 296058 274522 296146
rect 274630 296058 274810 296146
rect 275064 296058 275244 296146
rect 275352 296058 275532 296146
rect 275640 296058 275820 296146
rect 275928 296058 276108 296146
rect 276216 296058 276396 296146
rect 276504 296058 276684 296146
rect 276792 296058 276972 296146
rect 277080 296058 277260 296146
rect 277514 296058 277694 296146
rect 277802 296058 277982 296146
rect 278090 296058 278270 296146
rect 278378 296058 278558 296146
rect 278666 296058 278846 296146
rect 278954 296058 279134 296146
rect 279242 296058 279422 296146
rect 279530 296058 279710 296146
rect 279964 296058 280144 296146
rect 280252 296058 280432 296146
rect 280540 296058 280720 296146
rect 280828 296058 281008 296146
rect 281116 296058 281296 296146
rect 281404 296058 281584 296146
rect 281692 296058 281872 296146
rect 281980 296058 282160 296146
rect 282414 296058 282594 296146
rect 282702 296058 282882 296146
rect 282990 296058 283170 296146
rect 283278 296058 283458 296146
rect 283566 296058 283746 296146
rect 283854 296058 284034 296146
rect 284142 296058 284322 296146
rect 284430 296058 284610 296146
rect 284864 296058 285044 296146
rect 285152 296058 285332 296146
rect 285440 296058 285620 296146
rect 285728 296058 285908 296146
rect 286016 296058 286196 296146
rect 286304 296058 286484 296146
rect 286592 296058 286772 296146
rect 286880 296058 287060 296146
rect 287314 296058 287494 296146
rect 287602 296058 287782 296146
rect 287890 296058 288070 296146
rect 288178 296058 288358 296146
rect 288466 296058 288646 296146
rect 288754 296058 288934 296146
rect 289042 296058 289222 296146
rect 289330 296058 289510 296146
rect 289764 296058 289944 296146
rect 290052 296058 290232 296146
rect 290340 296058 290520 296146
rect 290628 296058 290808 296146
rect 290916 296058 291096 296146
rect 291204 296058 291384 296146
rect 291492 296058 291672 296146
rect 291780 296058 291960 296146
rect 292214 296058 292394 296146
rect 292502 296058 292682 296146
rect 292790 296058 292970 296146
rect 293078 296058 293258 296146
rect 293366 296058 293546 296146
rect 293654 296058 293834 296146
rect 293942 296058 294122 296146
rect 294230 296058 294410 296146
rect 294664 296058 294844 296146
rect 294952 296058 295132 296146
rect 295240 296058 295420 296146
rect 295528 296058 295708 296146
rect 295816 296058 295996 296146
rect 296104 296058 296284 296146
rect 296392 296058 296572 296146
rect 296680 296058 296860 296146
rect 297114 296058 297294 296146
rect 297402 296058 297582 296146
rect 297690 296058 297870 296146
rect 297978 296058 298158 296146
rect 298266 296058 298446 296146
rect 298554 296058 298734 296146
rect 298842 296058 299022 296146
rect 299130 296058 299310 296146
rect 299564 296058 299744 296146
rect 299852 296058 300032 296146
rect 300140 296058 300320 296146
rect 300428 296058 300608 296146
rect 300716 296058 300896 296146
rect 301004 296058 301184 296146
rect 301292 296058 301472 296146
rect 301580 296058 301760 296146
rect 302014 296058 302194 296146
rect 302302 296058 302482 296146
rect 302590 296058 302770 296146
rect 302878 296058 303058 296146
rect 303166 296058 303346 296146
rect 303454 296058 303634 296146
rect 303742 296058 303922 296146
rect 304030 296058 304210 296146
rect 304464 296058 304644 296146
rect 304752 296058 304932 296146
rect 305040 296058 305220 296146
rect 305328 296058 305508 296146
rect 305616 296058 305796 296146
rect 305904 296058 306084 296146
rect 306192 296058 306372 296146
rect 306480 296058 306660 296146
rect 306914 296058 307094 296146
rect 307202 296058 307382 296146
rect 307490 296058 307670 296146
rect 307778 296058 307958 296146
rect 308066 296058 308246 296146
rect 308354 296058 308534 296146
rect 308642 296058 308822 296146
rect 308930 296058 309110 296146
rect 309364 296058 309544 296146
rect 309652 296058 309832 296146
rect 309940 296058 310120 296146
rect 310228 296058 310408 296146
rect 310516 296058 310696 296146
rect 310804 296058 310984 296146
rect 311092 296058 311272 296146
rect 311380 296058 311560 296146
rect 311814 296058 311994 296146
rect 312102 296058 312282 296146
rect 312390 296058 312570 296146
rect 312678 296058 312858 296146
rect 312966 296058 313146 296146
rect 313254 296058 313434 296146
rect 313542 296058 313722 296146
rect 313830 296058 314010 296146
rect 314264 296058 314444 296146
rect 314552 296058 314732 296146
rect 314840 296058 315020 296146
rect 315128 296058 315308 296146
rect 315416 296058 315596 296146
rect 315704 296058 315884 296146
rect 315992 296058 316172 296146
rect 316280 296058 316460 296146
rect 316714 296058 316894 296146
rect 317002 296058 317182 296146
rect 317290 296058 317470 296146
rect 317578 296058 317758 296146
rect 317866 296058 318046 296146
rect 318154 296058 318334 296146
rect 318442 296058 318622 296146
rect 318730 296058 318910 296146
rect 319164 296058 319344 296146
rect 319452 296058 319632 296146
rect 319740 296058 319920 296146
rect 320028 296058 320208 296146
rect 320316 296058 320496 296146
rect 320604 296058 320784 296146
rect 320892 296058 321072 296146
rect 321180 296058 321360 296146
rect 321614 296058 321794 296146
rect 321902 296058 322082 296146
rect 322190 296058 322370 296146
rect 322478 296058 322658 296146
rect 322766 296058 322946 296146
rect 323054 296058 323234 296146
rect 323342 296058 323522 296146
rect 323630 296058 323810 296146
rect 324064 296058 324244 296146
rect 324352 296058 324532 296146
rect 324640 296058 324820 296146
rect 324928 296058 325108 296146
rect 325216 296058 325396 296146
rect 325504 296058 325684 296146
rect 325792 296058 325972 296146
rect 326080 296058 326260 296146
rect 326514 296058 326694 296146
rect 326802 296058 326982 296146
rect 327090 296058 327270 296146
rect 327378 296058 327558 296146
rect 327666 296058 327846 296146
rect 327954 296058 328134 296146
rect 328242 296058 328422 296146
rect 328530 296058 328710 296146
rect 328964 296058 329144 296146
rect 329252 296058 329432 296146
rect 329540 296058 329720 296146
rect 329828 296058 330008 296146
rect 330116 296058 330296 296146
rect 330404 296058 330584 296146
rect 330692 296058 330872 296146
rect 330980 296058 331160 296146
rect 331414 296058 331594 296146
rect 331702 296058 331882 296146
rect 331990 296058 332170 296146
rect 332278 296058 332458 296146
rect 332566 296058 332746 296146
rect 332854 296058 333034 296146
rect 333142 296058 333322 296146
rect 333430 296058 333610 296146
rect 333864 296058 334044 296146
rect 334152 296058 334332 296146
rect 334440 296058 334620 296146
rect 334728 296058 334908 296146
rect 335016 296058 335196 296146
rect 335304 296058 335484 296146
rect 335592 296058 335772 296146
rect 335880 296058 336060 296146
rect 336314 296058 336494 296146
rect 336602 296058 336782 296146
rect 336890 296058 337070 296146
rect 337178 296058 337358 296146
rect 337466 296058 337646 296146
rect 337754 296058 337934 296146
rect 338042 296058 338222 296146
rect 338330 296058 338510 296146
rect 338764 296058 338944 296146
rect 339052 296058 339232 296146
rect 339340 296058 339520 296146
rect 339628 296058 339808 296146
rect 339916 296058 340096 296146
rect 340204 296058 340384 296146
rect 340492 296058 340672 296146
rect 340780 296058 340960 296146
rect 341214 296058 341394 296146
rect 341502 296058 341682 296146
rect 341790 296058 341970 296146
rect 342078 296058 342258 296146
rect 342366 296058 342546 296146
rect 342654 296058 342834 296146
rect 342942 296058 343122 296146
rect 343230 296058 343410 296146
rect 343664 296058 343844 296146
rect 343952 296058 344132 296146
rect 344240 296058 344420 296146
rect 344528 296058 344708 296146
rect 344816 296058 344996 296146
rect 345104 296058 345284 296146
rect 345392 296058 345572 296146
rect 345680 296058 345860 296146
rect 346114 296058 346294 296146
rect 346402 296058 346582 296146
rect 346690 296058 346870 296146
rect 346978 296058 347158 296146
rect 347266 296058 347446 296146
rect 347554 296058 347734 296146
rect 347842 296058 348022 296146
rect 348130 296058 348310 296146
rect 348564 296058 348744 296146
rect 348852 296058 349032 296146
rect 349140 296058 349320 296146
rect 349428 296058 349608 296146
rect 349716 296058 349896 296146
rect 350004 296058 350184 296146
rect 350292 296058 350472 296146
rect 350580 296058 350760 296146
rect 351014 296058 351194 296146
rect 351302 296058 351482 296146
rect 351590 296058 351770 296146
rect 351878 296058 352058 296146
rect 352166 296058 352346 296146
rect 352454 296058 352634 296146
rect 352742 296058 352922 296146
rect 353030 296058 353210 296146
rect 353464 296058 353644 296146
rect 353752 296058 353932 296146
rect 354040 296058 354220 296146
rect 354328 296058 354508 296146
rect 354616 296058 354796 296146
rect 354904 296058 355084 296146
rect 355192 296058 355372 296146
rect 355480 296058 355660 296146
rect 355914 296058 356094 296146
rect 356202 296058 356382 296146
rect 356490 296058 356670 296146
rect 356778 296058 356958 296146
rect 357066 296058 357246 296146
rect 357354 296058 357534 296146
rect 357642 296058 357822 296146
rect 357930 296058 358110 296146
rect 358364 296058 358544 296146
rect 358652 296058 358832 296146
rect 358940 296058 359120 296146
rect 359228 296058 359408 296146
rect 359516 296058 359696 296146
rect 359804 296058 359984 296146
rect 360092 296058 360272 296146
rect 360380 296058 360560 296146
rect 360814 296058 360994 296146
rect 361102 296058 361282 296146
rect 361390 296058 361570 296146
rect 361678 296058 361858 296146
rect 361966 296058 362146 296146
rect 362254 296058 362434 296146
rect 362542 296058 362722 296146
rect 362830 296058 363010 296146
rect 363264 296058 363444 296146
rect 363552 296058 363732 296146
rect 363840 296058 364020 296146
rect 364128 296058 364308 296146
rect 364416 296058 364596 296146
rect 364704 296058 364884 296146
rect 364992 296058 365172 296146
rect 365280 296058 365460 296146
rect 365714 296058 365894 296146
rect 366002 296058 366182 296146
rect 366290 296058 366470 296146
rect 366578 296058 366758 296146
rect 366866 296058 367046 296146
rect 367154 296058 367334 296146
rect 367442 296058 367622 296146
rect 367730 296058 367910 296146
rect 243214 295582 243394 295670
rect 243502 295582 243682 295670
rect 243790 295582 243970 295670
rect 244078 295582 244258 295670
rect 244366 295582 244546 295670
rect 244654 295582 244834 295670
rect 244942 295582 245122 295670
rect 245230 295582 245410 295670
rect 245664 295582 245844 295670
rect 245952 295582 246132 295670
rect 246240 295582 246420 295670
rect 246528 295582 246708 295670
rect 246816 295582 246996 295670
rect 247104 295582 247284 295670
rect 247392 295582 247572 295670
rect 247680 295582 247860 295670
rect 248114 295582 248294 295670
rect 248402 295582 248582 295670
rect 248690 295582 248870 295670
rect 248978 295582 249158 295670
rect 249266 295582 249446 295670
rect 249554 295582 249734 295670
rect 249842 295582 250022 295670
rect 250130 295582 250310 295670
rect 250564 295582 250744 295670
rect 250852 295582 251032 295670
rect 251140 295582 251320 295670
rect 251428 295582 251608 295670
rect 251716 295582 251896 295670
rect 252004 295582 252184 295670
rect 252292 295582 252472 295670
rect 252580 295582 252760 295670
rect 253014 295582 253194 295670
rect 253302 295582 253482 295670
rect 253590 295582 253770 295670
rect 253878 295582 254058 295670
rect 254166 295582 254346 295670
rect 254454 295582 254634 295670
rect 254742 295582 254922 295670
rect 255030 295582 255210 295670
rect 255464 295582 255644 295670
rect 255752 295582 255932 295670
rect 256040 295582 256220 295670
rect 256328 295582 256508 295670
rect 256616 295582 256796 295670
rect 256904 295582 257084 295670
rect 257192 295582 257372 295670
rect 257480 295582 257660 295670
rect 257914 295582 258094 295670
rect 258202 295582 258382 295670
rect 258490 295582 258670 295670
rect 258778 295582 258958 295670
rect 259066 295582 259246 295670
rect 259354 295582 259534 295670
rect 259642 295582 259822 295670
rect 259930 295582 260110 295670
rect 260364 295582 260544 295670
rect 260652 295582 260832 295670
rect 260940 295582 261120 295670
rect 261228 295582 261408 295670
rect 261516 295582 261696 295670
rect 261804 295582 261984 295670
rect 262092 295582 262272 295670
rect 262380 295582 262560 295670
rect 262814 295582 262994 295670
rect 263102 295582 263282 295670
rect 263390 295582 263570 295670
rect 263678 295582 263858 295670
rect 263966 295582 264146 295670
rect 264254 295582 264434 295670
rect 264542 295582 264722 295670
rect 264830 295582 265010 295670
rect 265264 295582 265444 295670
rect 265552 295582 265732 295670
rect 265840 295582 266020 295670
rect 266128 295582 266308 295670
rect 266416 295582 266596 295670
rect 266704 295582 266884 295670
rect 266992 295582 267172 295670
rect 267280 295582 267460 295670
rect 267714 295582 267894 295670
rect 268002 295582 268182 295670
rect 268290 295582 268470 295670
rect 268578 295582 268758 295670
rect 268866 295582 269046 295670
rect 269154 295582 269334 295670
rect 269442 295582 269622 295670
rect 269730 295582 269910 295670
rect 270164 295582 270344 295670
rect 270452 295582 270632 295670
rect 270740 295582 270920 295670
rect 271028 295582 271208 295670
rect 271316 295582 271496 295670
rect 271604 295582 271784 295670
rect 271892 295582 272072 295670
rect 272180 295582 272360 295670
rect 272614 295582 272794 295670
rect 272902 295582 273082 295670
rect 273190 295582 273370 295670
rect 273478 295582 273658 295670
rect 273766 295582 273946 295670
rect 274054 295582 274234 295670
rect 274342 295582 274522 295670
rect 274630 295582 274810 295670
rect 275064 295582 275244 295670
rect 275352 295582 275532 295670
rect 275640 295582 275820 295670
rect 275928 295582 276108 295670
rect 276216 295582 276396 295670
rect 276504 295582 276684 295670
rect 276792 295582 276972 295670
rect 277080 295582 277260 295670
rect 277514 295582 277694 295670
rect 277802 295582 277982 295670
rect 278090 295582 278270 295670
rect 278378 295582 278558 295670
rect 278666 295582 278846 295670
rect 278954 295582 279134 295670
rect 279242 295582 279422 295670
rect 279530 295582 279710 295670
rect 279964 295582 280144 295670
rect 280252 295582 280432 295670
rect 280540 295582 280720 295670
rect 280828 295582 281008 295670
rect 281116 295582 281296 295670
rect 281404 295582 281584 295670
rect 281692 295582 281872 295670
rect 281980 295582 282160 295670
rect 282414 295582 282594 295670
rect 282702 295582 282882 295670
rect 282990 295582 283170 295670
rect 283278 295582 283458 295670
rect 283566 295582 283746 295670
rect 283854 295582 284034 295670
rect 284142 295582 284322 295670
rect 284430 295582 284610 295670
rect 284864 295582 285044 295670
rect 285152 295582 285332 295670
rect 285440 295582 285620 295670
rect 285728 295582 285908 295670
rect 286016 295582 286196 295670
rect 286304 295582 286484 295670
rect 286592 295582 286772 295670
rect 286880 295582 287060 295670
rect 287314 295582 287494 295670
rect 287602 295582 287782 295670
rect 287890 295582 288070 295670
rect 288178 295582 288358 295670
rect 288466 295582 288646 295670
rect 288754 295582 288934 295670
rect 289042 295582 289222 295670
rect 289330 295582 289510 295670
rect 289764 295582 289944 295670
rect 290052 295582 290232 295670
rect 290340 295582 290520 295670
rect 290628 295582 290808 295670
rect 290916 295582 291096 295670
rect 291204 295582 291384 295670
rect 291492 295582 291672 295670
rect 291780 295582 291960 295670
rect 292214 295582 292394 295670
rect 292502 295582 292682 295670
rect 292790 295582 292970 295670
rect 293078 295582 293258 295670
rect 293366 295582 293546 295670
rect 293654 295582 293834 295670
rect 293942 295582 294122 295670
rect 294230 295582 294410 295670
rect 294664 295582 294844 295670
rect 294952 295582 295132 295670
rect 295240 295582 295420 295670
rect 295528 295582 295708 295670
rect 295816 295582 295996 295670
rect 296104 295582 296284 295670
rect 296392 295582 296572 295670
rect 296680 295582 296860 295670
rect 297114 295582 297294 295670
rect 297402 295582 297582 295670
rect 297690 295582 297870 295670
rect 297978 295582 298158 295670
rect 298266 295582 298446 295670
rect 298554 295582 298734 295670
rect 298842 295582 299022 295670
rect 299130 295582 299310 295670
rect 299564 295582 299744 295670
rect 299852 295582 300032 295670
rect 300140 295582 300320 295670
rect 300428 295582 300608 295670
rect 300716 295582 300896 295670
rect 301004 295582 301184 295670
rect 301292 295582 301472 295670
rect 301580 295582 301760 295670
rect 302014 295582 302194 295670
rect 302302 295582 302482 295670
rect 302590 295582 302770 295670
rect 302878 295582 303058 295670
rect 303166 295582 303346 295670
rect 303454 295582 303634 295670
rect 303742 295582 303922 295670
rect 304030 295582 304210 295670
rect 304464 295582 304644 295670
rect 304752 295582 304932 295670
rect 305040 295582 305220 295670
rect 305328 295582 305508 295670
rect 305616 295582 305796 295670
rect 305904 295582 306084 295670
rect 306192 295582 306372 295670
rect 306480 295582 306660 295670
rect 306914 295582 307094 295670
rect 307202 295582 307382 295670
rect 307490 295582 307670 295670
rect 307778 295582 307958 295670
rect 308066 295582 308246 295670
rect 308354 295582 308534 295670
rect 308642 295582 308822 295670
rect 308930 295582 309110 295670
rect 309364 295582 309544 295670
rect 309652 295582 309832 295670
rect 309940 295582 310120 295670
rect 310228 295582 310408 295670
rect 310516 295582 310696 295670
rect 310804 295582 310984 295670
rect 311092 295582 311272 295670
rect 311380 295582 311560 295670
rect 311814 295582 311994 295670
rect 312102 295582 312282 295670
rect 312390 295582 312570 295670
rect 312678 295582 312858 295670
rect 312966 295582 313146 295670
rect 313254 295582 313434 295670
rect 313542 295582 313722 295670
rect 313830 295582 314010 295670
rect 314264 295582 314444 295670
rect 314552 295582 314732 295670
rect 314840 295582 315020 295670
rect 315128 295582 315308 295670
rect 315416 295582 315596 295670
rect 315704 295582 315884 295670
rect 315992 295582 316172 295670
rect 316280 295582 316460 295670
rect 316714 295582 316894 295670
rect 317002 295582 317182 295670
rect 317290 295582 317470 295670
rect 317578 295582 317758 295670
rect 317866 295582 318046 295670
rect 318154 295582 318334 295670
rect 318442 295582 318622 295670
rect 318730 295582 318910 295670
rect 319164 295582 319344 295670
rect 319452 295582 319632 295670
rect 319740 295582 319920 295670
rect 320028 295582 320208 295670
rect 320316 295582 320496 295670
rect 320604 295582 320784 295670
rect 320892 295582 321072 295670
rect 321180 295582 321360 295670
rect 321614 295582 321794 295670
rect 321902 295582 322082 295670
rect 322190 295582 322370 295670
rect 322478 295582 322658 295670
rect 322766 295582 322946 295670
rect 323054 295582 323234 295670
rect 323342 295582 323522 295670
rect 323630 295582 323810 295670
rect 324064 295582 324244 295670
rect 324352 295582 324532 295670
rect 324640 295582 324820 295670
rect 324928 295582 325108 295670
rect 325216 295582 325396 295670
rect 325504 295582 325684 295670
rect 325792 295582 325972 295670
rect 326080 295582 326260 295670
rect 326514 295582 326694 295670
rect 326802 295582 326982 295670
rect 327090 295582 327270 295670
rect 327378 295582 327558 295670
rect 327666 295582 327846 295670
rect 327954 295582 328134 295670
rect 328242 295582 328422 295670
rect 328530 295582 328710 295670
rect 328964 295582 329144 295670
rect 329252 295582 329432 295670
rect 329540 295582 329720 295670
rect 329828 295582 330008 295670
rect 330116 295582 330296 295670
rect 330404 295582 330584 295670
rect 330692 295582 330872 295670
rect 330980 295582 331160 295670
rect 331414 295582 331594 295670
rect 331702 295582 331882 295670
rect 331990 295582 332170 295670
rect 332278 295582 332458 295670
rect 332566 295582 332746 295670
rect 332854 295582 333034 295670
rect 333142 295582 333322 295670
rect 333430 295582 333610 295670
rect 333864 295582 334044 295670
rect 334152 295582 334332 295670
rect 334440 295582 334620 295670
rect 334728 295582 334908 295670
rect 335016 295582 335196 295670
rect 335304 295582 335484 295670
rect 335592 295582 335772 295670
rect 335880 295582 336060 295670
rect 336314 295582 336494 295670
rect 336602 295582 336782 295670
rect 336890 295582 337070 295670
rect 337178 295582 337358 295670
rect 337466 295582 337646 295670
rect 337754 295582 337934 295670
rect 338042 295582 338222 295670
rect 338330 295582 338510 295670
rect 338764 295582 338944 295670
rect 339052 295582 339232 295670
rect 339340 295582 339520 295670
rect 339628 295582 339808 295670
rect 339916 295582 340096 295670
rect 340204 295582 340384 295670
rect 340492 295582 340672 295670
rect 340780 295582 340960 295670
rect 341214 295582 341394 295670
rect 341502 295582 341682 295670
rect 341790 295582 341970 295670
rect 342078 295582 342258 295670
rect 342366 295582 342546 295670
rect 342654 295582 342834 295670
rect 342942 295582 343122 295670
rect 343230 295582 343410 295670
rect 343664 295582 343844 295670
rect 343952 295582 344132 295670
rect 344240 295582 344420 295670
rect 344528 295582 344708 295670
rect 344816 295582 344996 295670
rect 345104 295582 345284 295670
rect 345392 295582 345572 295670
rect 345680 295582 345860 295670
rect 346114 295582 346294 295670
rect 346402 295582 346582 295670
rect 346690 295582 346870 295670
rect 346978 295582 347158 295670
rect 347266 295582 347446 295670
rect 347554 295582 347734 295670
rect 347842 295582 348022 295670
rect 348130 295582 348310 295670
rect 348564 295582 348744 295670
rect 348852 295582 349032 295670
rect 349140 295582 349320 295670
rect 349428 295582 349608 295670
rect 349716 295582 349896 295670
rect 350004 295582 350184 295670
rect 350292 295582 350472 295670
rect 350580 295582 350760 295670
rect 351014 295582 351194 295670
rect 351302 295582 351482 295670
rect 351590 295582 351770 295670
rect 351878 295582 352058 295670
rect 352166 295582 352346 295670
rect 352454 295582 352634 295670
rect 352742 295582 352922 295670
rect 353030 295582 353210 295670
rect 353464 295582 353644 295670
rect 353752 295582 353932 295670
rect 354040 295582 354220 295670
rect 354328 295582 354508 295670
rect 354616 295582 354796 295670
rect 354904 295582 355084 295670
rect 355192 295582 355372 295670
rect 355480 295582 355660 295670
rect 355914 295582 356094 295670
rect 356202 295582 356382 295670
rect 356490 295582 356670 295670
rect 356778 295582 356958 295670
rect 357066 295582 357246 295670
rect 357354 295582 357534 295670
rect 357642 295582 357822 295670
rect 357930 295582 358110 295670
rect 358364 295582 358544 295670
rect 358652 295582 358832 295670
rect 358940 295582 359120 295670
rect 359228 295582 359408 295670
rect 359516 295582 359696 295670
rect 359804 295582 359984 295670
rect 360092 295582 360272 295670
rect 360380 295582 360560 295670
rect 360814 295582 360994 295670
rect 361102 295582 361282 295670
rect 361390 295582 361570 295670
rect 361678 295582 361858 295670
rect 361966 295582 362146 295670
rect 362254 295582 362434 295670
rect 362542 295582 362722 295670
rect 362830 295582 363010 295670
rect 363264 295582 363444 295670
rect 363552 295582 363732 295670
rect 363840 295582 364020 295670
rect 364128 295582 364308 295670
rect 364416 295582 364596 295670
rect 364704 295582 364884 295670
rect 364992 295582 365172 295670
rect 365280 295582 365460 295670
rect 365714 295582 365894 295670
rect 366002 295582 366182 295670
rect 366290 295582 366470 295670
rect 366578 295582 366758 295670
rect 366866 295582 367046 295670
rect 367154 295582 367334 295670
rect 367442 295582 367622 295670
rect 367730 295582 367910 295670
rect 243214 295366 243394 295454
rect 243502 295366 243682 295454
rect 243790 295366 243970 295454
rect 244078 295366 244258 295454
rect 244366 295366 244546 295454
rect 244654 295366 244834 295454
rect 244942 295366 245122 295454
rect 245230 295366 245410 295454
rect 245664 295366 245844 295454
rect 245952 295366 246132 295454
rect 246240 295366 246420 295454
rect 246528 295366 246708 295454
rect 246816 295366 246996 295454
rect 247104 295366 247284 295454
rect 247392 295366 247572 295454
rect 247680 295366 247860 295454
rect 248114 295366 248294 295454
rect 248402 295366 248582 295454
rect 248690 295366 248870 295454
rect 248978 295366 249158 295454
rect 249266 295366 249446 295454
rect 249554 295366 249734 295454
rect 249842 295366 250022 295454
rect 250130 295366 250310 295454
rect 250564 295366 250744 295454
rect 250852 295366 251032 295454
rect 251140 295366 251320 295454
rect 251428 295366 251608 295454
rect 251716 295366 251896 295454
rect 252004 295366 252184 295454
rect 252292 295366 252472 295454
rect 252580 295366 252760 295454
rect 253014 295366 253194 295454
rect 253302 295366 253482 295454
rect 253590 295366 253770 295454
rect 253878 295366 254058 295454
rect 254166 295366 254346 295454
rect 254454 295366 254634 295454
rect 254742 295366 254922 295454
rect 255030 295366 255210 295454
rect 255464 295366 255644 295454
rect 255752 295366 255932 295454
rect 256040 295366 256220 295454
rect 256328 295366 256508 295454
rect 256616 295366 256796 295454
rect 256904 295366 257084 295454
rect 257192 295366 257372 295454
rect 257480 295366 257660 295454
rect 257914 295366 258094 295454
rect 258202 295366 258382 295454
rect 258490 295366 258670 295454
rect 258778 295366 258958 295454
rect 259066 295366 259246 295454
rect 259354 295366 259534 295454
rect 259642 295366 259822 295454
rect 259930 295366 260110 295454
rect 260364 295366 260544 295454
rect 260652 295366 260832 295454
rect 260940 295366 261120 295454
rect 261228 295366 261408 295454
rect 261516 295366 261696 295454
rect 261804 295366 261984 295454
rect 262092 295366 262272 295454
rect 262380 295366 262560 295454
rect 262814 295366 262994 295454
rect 263102 295366 263282 295454
rect 263390 295366 263570 295454
rect 263678 295366 263858 295454
rect 263966 295366 264146 295454
rect 264254 295366 264434 295454
rect 264542 295366 264722 295454
rect 264830 295366 265010 295454
rect 265264 295366 265444 295454
rect 265552 295366 265732 295454
rect 265840 295366 266020 295454
rect 266128 295366 266308 295454
rect 266416 295366 266596 295454
rect 266704 295366 266884 295454
rect 266992 295366 267172 295454
rect 267280 295366 267460 295454
rect 267714 295366 267894 295454
rect 268002 295366 268182 295454
rect 268290 295366 268470 295454
rect 268578 295366 268758 295454
rect 268866 295366 269046 295454
rect 269154 295366 269334 295454
rect 269442 295366 269622 295454
rect 269730 295366 269910 295454
rect 270164 295366 270344 295454
rect 270452 295366 270632 295454
rect 270740 295366 270920 295454
rect 271028 295366 271208 295454
rect 271316 295366 271496 295454
rect 271604 295366 271784 295454
rect 271892 295366 272072 295454
rect 272180 295366 272360 295454
rect 272614 295366 272794 295454
rect 272902 295366 273082 295454
rect 273190 295366 273370 295454
rect 273478 295366 273658 295454
rect 273766 295366 273946 295454
rect 274054 295366 274234 295454
rect 274342 295366 274522 295454
rect 274630 295366 274810 295454
rect 275064 295366 275244 295454
rect 275352 295366 275532 295454
rect 275640 295366 275820 295454
rect 275928 295366 276108 295454
rect 276216 295366 276396 295454
rect 276504 295366 276684 295454
rect 276792 295366 276972 295454
rect 277080 295366 277260 295454
rect 277514 295366 277694 295454
rect 277802 295366 277982 295454
rect 278090 295366 278270 295454
rect 278378 295366 278558 295454
rect 278666 295366 278846 295454
rect 278954 295366 279134 295454
rect 279242 295366 279422 295454
rect 279530 295366 279710 295454
rect 279964 295366 280144 295454
rect 280252 295366 280432 295454
rect 280540 295366 280720 295454
rect 280828 295366 281008 295454
rect 281116 295366 281296 295454
rect 281404 295366 281584 295454
rect 281692 295366 281872 295454
rect 281980 295366 282160 295454
rect 282414 295366 282594 295454
rect 282702 295366 282882 295454
rect 282990 295366 283170 295454
rect 283278 295366 283458 295454
rect 283566 295366 283746 295454
rect 283854 295366 284034 295454
rect 284142 295366 284322 295454
rect 284430 295366 284610 295454
rect 284864 295366 285044 295454
rect 285152 295366 285332 295454
rect 285440 295366 285620 295454
rect 285728 295366 285908 295454
rect 286016 295366 286196 295454
rect 286304 295366 286484 295454
rect 286592 295366 286772 295454
rect 286880 295366 287060 295454
rect 287314 295366 287494 295454
rect 287602 295366 287782 295454
rect 287890 295366 288070 295454
rect 288178 295366 288358 295454
rect 288466 295366 288646 295454
rect 288754 295366 288934 295454
rect 289042 295366 289222 295454
rect 289330 295366 289510 295454
rect 289764 295366 289944 295454
rect 290052 295366 290232 295454
rect 290340 295366 290520 295454
rect 290628 295366 290808 295454
rect 290916 295366 291096 295454
rect 291204 295366 291384 295454
rect 291492 295366 291672 295454
rect 291780 295366 291960 295454
rect 292214 295366 292394 295454
rect 292502 295366 292682 295454
rect 292790 295366 292970 295454
rect 293078 295366 293258 295454
rect 293366 295366 293546 295454
rect 293654 295366 293834 295454
rect 293942 295366 294122 295454
rect 294230 295366 294410 295454
rect 294664 295366 294844 295454
rect 294952 295366 295132 295454
rect 295240 295366 295420 295454
rect 295528 295366 295708 295454
rect 295816 295366 295996 295454
rect 296104 295366 296284 295454
rect 296392 295366 296572 295454
rect 296680 295366 296860 295454
rect 297114 295366 297294 295454
rect 297402 295366 297582 295454
rect 297690 295366 297870 295454
rect 297978 295366 298158 295454
rect 298266 295366 298446 295454
rect 298554 295366 298734 295454
rect 298842 295366 299022 295454
rect 299130 295366 299310 295454
rect 299564 295366 299744 295454
rect 299852 295366 300032 295454
rect 300140 295366 300320 295454
rect 300428 295366 300608 295454
rect 300716 295366 300896 295454
rect 301004 295366 301184 295454
rect 301292 295366 301472 295454
rect 301580 295366 301760 295454
rect 302014 295366 302194 295454
rect 302302 295366 302482 295454
rect 302590 295366 302770 295454
rect 302878 295366 303058 295454
rect 303166 295366 303346 295454
rect 303454 295366 303634 295454
rect 303742 295366 303922 295454
rect 304030 295366 304210 295454
rect 304464 295366 304644 295454
rect 304752 295366 304932 295454
rect 305040 295366 305220 295454
rect 305328 295366 305508 295454
rect 305616 295366 305796 295454
rect 305904 295366 306084 295454
rect 306192 295366 306372 295454
rect 306480 295366 306660 295454
rect 306914 295366 307094 295454
rect 307202 295366 307382 295454
rect 307490 295366 307670 295454
rect 307778 295366 307958 295454
rect 308066 295366 308246 295454
rect 308354 295366 308534 295454
rect 308642 295366 308822 295454
rect 308930 295366 309110 295454
rect 309364 295366 309544 295454
rect 309652 295366 309832 295454
rect 309940 295366 310120 295454
rect 310228 295366 310408 295454
rect 310516 295366 310696 295454
rect 310804 295366 310984 295454
rect 311092 295366 311272 295454
rect 311380 295366 311560 295454
rect 311814 295366 311994 295454
rect 312102 295366 312282 295454
rect 312390 295366 312570 295454
rect 312678 295366 312858 295454
rect 312966 295366 313146 295454
rect 313254 295366 313434 295454
rect 313542 295366 313722 295454
rect 313830 295366 314010 295454
rect 314264 295366 314444 295454
rect 314552 295366 314732 295454
rect 314840 295366 315020 295454
rect 315128 295366 315308 295454
rect 315416 295366 315596 295454
rect 315704 295366 315884 295454
rect 315992 295366 316172 295454
rect 316280 295366 316460 295454
rect 316714 295366 316894 295454
rect 317002 295366 317182 295454
rect 317290 295366 317470 295454
rect 317578 295366 317758 295454
rect 317866 295366 318046 295454
rect 318154 295366 318334 295454
rect 318442 295366 318622 295454
rect 318730 295366 318910 295454
rect 319164 295366 319344 295454
rect 319452 295366 319632 295454
rect 319740 295366 319920 295454
rect 320028 295366 320208 295454
rect 320316 295366 320496 295454
rect 320604 295366 320784 295454
rect 320892 295366 321072 295454
rect 321180 295366 321360 295454
rect 321614 295366 321794 295454
rect 321902 295366 322082 295454
rect 322190 295366 322370 295454
rect 322478 295366 322658 295454
rect 322766 295366 322946 295454
rect 323054 295366 323234 295454
rect 323342 295366 323522 295454
rect 323630 295366 323810 295454
rect 324064 295366 324244 295454
rect 324352 295366 324532 295454
rect 324640 295366 324820 295454
rect 324928 295366 325108 295454
rect 325216 295366 325396 295454
rect 325504 295366 325684 295454
rect 325792 295366 325972 295454
rect 326080 295366 326260 295454
rect 326514 295366 326694 295454
rect 326802 295366 326982 295454
rect 327090 295366 327270 295454
rect 327378 295366 327558 295454
rect 327666 295366 327846 295454
rect 327954 295366 328134 295454
rect 328242 295366 328422 295454
rect 328530 295366 328710 295454
rect 328964 295366 329144 295454
rect 329252 295366 329432 295454
rect 329540 295366 329720 295454
rect 329828 295366 330008 295454
rect 330116 295366 330296 295454
rect 330404 295366 330584 295454
rect 330692 295366 330872 295454
rect 330980 295366 331160 295454
rect 331414 295366 331594 295454
rect 331702 295366 331882 295454
rect 331990 295366 332170 295454
rect 332278 295366 332458 295454
rect 332566 295366 332746 295454
rect 332854 295366 333034 295454
rect 333142 295366 333322 295454
rect 333430 295366 333610 295454
rect 333864 295366 334044 295454
rect 334152 295366 334332 295454
rect 334440 295366 334620 295454
rect 334728 295366 334908 295454
rect 335016 295366 335196 295454
rect 335304 295366 335484 295454
rect 335592 295366 335772 295454
rect 335880 295366 336060 295454
rect 336314 295366 336494 295454
rect 336602 295366 336782 295454
rect 336890 295366 337070 295454
rect 337178 295366 337358 295454
rect 337466 295366 337646 295454
rect 337754 295366 337934 295454
rect 338042 295366 338222 295454
rect 338330 295366 338510 295454
rect 338764 295366 338944 295454
rect 339052 295366 339232 295454
rect 339340 295366 339520 295454
rect 339628 295366 339808 295454
rect 339916 295366 340096 295454
rect 340204 295366 340384 295454
rect 340492 295366 340672 295454
rect 340780 295366 340960 295454
rect 341214 295366 341394 295454
rect 341502 295366 341682 295454
rect 341790 295366 341970 295454
rect 342078 295366 342258 295454
rect 342366 295366 342546 295454
rect 342654 295366 342834 295454
rect 342942 295366 343122 295454
rect 343230 295366 343410 295454
rect 343664 295366 343844 295454
rect 343952 295366 344132 295454
rect 344240 295366 344420 295454
rect 344528 295366 344708 295454
rect 344816 295366 344996 295454
rect 345104 295366 345284 295454
rect 345392 295366 345572 295454
rect 345680 295366 345860 295454
rect 346114 295366 346294 295454
rect 346402 295366 346582 295454
rect 346690 295366 346870 295454
rect 346978 295366 347158 295454
rect 347266 295366 347446 295454
rect 347554 295366 347734 295454
rect 347842 295366 348022 295454
rect 348130 295366 348310 295454
rect 348564 295366 348744 295454
rect 348852 295366 349032 295454
rect 349140 295366 349320 295454
rect 349428 295366 349608 295454
rect 349716 295366 349896 295454
rect 350004 295366 350184 295454
rect 350292 295366 350472 295454
rect 350580 295366 350760 295454
rect 351014 295366 351194 295454
rect 351302 295366 351482 295454
rect 351590 295366 351770 295454
rect 351878 295366 352058 295454
rect 352166 295366 352346 295454
rect 352454 295366 352634 295454
rect 352742 295366 352922 295454
rect 353030 295366 353210 295454
rect 353464 295366 353644 295454
rect 353752 295366 353932 295454
rect 354040 295366 354220 295454
rect 354328 295366 354508 295454
rect 354616 295366 354796 295454
rect 354904 295366 355084 295454
rect 355192 295366 355372 295454
rect 355480 295366 355660 295454
rect 355914 295366 356094 295454
rect 356202 295366 356382 295454
rect 356490 295366 356670 295454
rect 356778 295366 356958 295454
rect 357066 295366 357246 295454
rect 357354 295366 357534 295454
rect 357642 295366 357822 295454
rect 357930 295366 358110 295454
rect 358364 295366 358544 295454
rect 358652 295366 358832 295454
rect 358940 295366 359120 295454
rect 359228 295366 359408 295454
rect 359516 295366 359696 295454
rect 359804 295366 359984 295454
rect 360092 295366 360272 295454
rect 360380 295366 360560 295454
rect 360814 295366 360994 295454
rect 361102 295366 361282 295454
rect 361390 295366 361570 295454
rect 361678 295366 361858 295454
rect 361966 295366 362146 295454
rect 362254 295366 362434 295454
rect 362542 295366 362722 295454
rect 362830 295366 363010 295454
rect 363264 295366 363444 295454
rect 363552 295366 363732 295454
rect 363840 295366 364020 295454
rect 364128 295366 364308 295454
rect 364416 295366 364596 295454
rect 364704 295366 364884 295454
rect 364992 295366 365172 295454
rect 365280 295366 365460 295454
rect 365714 295366 365894 295454
rect 366002 295366 366182 295454
rect 366290 295366 366470 295454
rect 366578 295366 366758 295454
rect 366866 295366 367046 295454
rect 367154 295366 367334 295454
rect 367442 295366 367622 295454
rect 367730 295366 367910 295454
rect 243214 294890 243394 294978
rect 243502 294890 243682 294978
rect 243790 294890 243970 294978
rect 244078 294890 244258 294978
rect 244366 294890 244546 294978
rect 244654 294890 244834 294978
rect 244942 294890 245122 294978
rect 245230 294890 245410 294978
rect 245664 294890 245844 294978
rect 245952 294890 246132 294978
rect 246240 294890 246420 294978
rect 246528 294890 246708 294978
rect 246816 294890 246996 294978
rect 247104 294890 247284 294978
rect 247392 294890 247572 294978
rect 247680 294890 247860 294978
rect 248114 294890 248294 294978
rect 248402 294890 248582 294978
rect 248690 294890 248870 294978
rect 248978 294890 249158 294978
rect 249266 294890 249446 294978
rect 249554 294890 249734 294978
rect 249842 294890 250022 294978
rect 250130 294890 250310 294978
rect 250564 294890 250744 294978
rect 250852 294890 251032 294978
rect 251140 294890 251320 294978
rect 251428 294890 251608 294978
rect 251716 294890 251896 294978
rect 252004 294890 252184 294978
rect 252292 294890 252472 294978
rect 252580 294890 252760 294978
rect 253014 294890 253194 294978
rect 253302 294890 253482 294978
rect 253590 294890 253770 294978
rect 253878 294890 254058 294978
rect 254166 294890 254346 294978
rect 254454 294890 254634 294978
rect 254742 294890 254922 294978
rect 255030 294890 255210 294978
rect 255464 294890 255644 294978
rect 255752 294890 255932 294978
rect 256040 294890 256220 294978
rect 256328 294890 256508 294978
rect 256616 294890 256796 294978
rect 256904 294890 257084 294978
rect 257192 294890 257372 294978
rect 257480 294890 257660 294978
rect 257914 294890 258094 294978
rect 258202 294890 258382 294978
rect 258490 294890 258670 294978
rect 258778 294890 258958 294978
rect 259066 294890 259246 294978
rect 259354 294890 259534 294978
rect 259642 294890 259822 294978
rect 259930 294890 260110 294978
rect 260364 294890 260544 294978
rect 260652 294890 260832 294978
rect 260940 294890 261120 294978
rect 261228 294890 261408 294978
rect 261516 294890 261696 294978
rect 261804 294890 261984 294978
rect 262092 294890 262272 294978
rect 262380 294890 262560 294978
rect 262814 294890 262994 294978
rect 263102 294890 263282 294978
rect 263390 294890 263570 294978
rect 263678 294890 263858 294978
rect 263966 294890 264146 294978
rect 264254 294890 264434 294978
rect 264542 294890 264722 294978
rect 264830 294890 265010 294978
rect 265264 294890 265444 294978
rect 265552 294890 265732 294978
rect 265840 294890 266020 294978
rect 266128 294890 266308 294978
rect 266416 294890 266596 294978
rect 266704 294890 266884 294978
rect 266992 294890 267172 294978
rect 267280 294890 267460 294978
rect 267714 294890 267894 294978
rect 268002 294890 268182 294978
rect 268290 294890 268470 294978
rect 268578 294890 268758 294978
rect 268866 294890 269046 294978
rect 269154 294890 269334 294978
rect 269442 294890 269622 294978
rect 269730 294890 269910 294978
rect 270164 294890 270344 294978
rect 270452 294890 270632 294978
rect 270740 294890 270920 294978
rect 271028 294890 271208 294978
rect 271316 294890 271496 294978
rect 271604 294890 271784 294978
rect 271892 294890 272072 294978
rect 272180 294890 272360 294978
rect 272614 294890 272794 294978
rect 272902 294890 273082 294978
rect 273190 294890 273370 294978
rect 273478 294890 273658 294978
rect 273766 294890 273946 294978
rect 274054 294890 274234 294978
rect 274342 294890 274522 294978
rect 274630 294890 274810 294978
rect 275064 294890 275244 294978
rect 275352 294890 275532 294978
rect 275640 294890 275820 294978
rect 275928 294890 276108 294978
rect 276216 294890 276396 294978
rect 276504 294890 276684 294978
rect 276792 294890 276972 294978
rect 277080 294890 277260 294978
rect 277514 294890 277694 294978
rect 277802 294890 277982 294978
rect 278090 294890 278270 294978
rect 278378 294890 278558 294978
rect 278666 294890 278846 294978
rect 278954 294890 279134 294978
rect 279242 294890 279422 294978
rect 279530 294890 279710 294978
rect 279964 294890 280144 294978
rect 280252 294890 280432 294978
rect 280540 294890 280720 294978
rect 280828 294890 281008 294978
rect 281116 294890 281296 294978
rect 281404 294890 281584 294978
rect 281692 294890 281872 294978
rect 281980 294890 282160 294978
rect 282414 294890 282594 294978
rect 282702 294890 282882 294978
rect 282990 294890 283170 294978
rect 283278 294890 283458 294978
rect 283566 294890 283746 294978
rect 283854 294890 284034 294978
rect 284142 294890 284322 294978
rect 284430 294890 284610 294978
rect 284864 294890 285044 294978
rect 285152 294890 285332 294978
rect 285440 294890 285620 294978
rect 285728 294890 285908 294978
rect 286016 294890 286196 294978
rect 286304 294890 286484 294978
rect 286592 294890 286772 294978
rect 286880 294890 287060 294978
rect 287314 294890 287494 294978
rect 287602 294890 287782 294978
rect 287890 294890 288070 294978
rect 288178 294890 288358 294978
rect 288466 294890 288646 294978
rect 288754 294890 288934 294978
rect 289042 294890 289222 294978
rect 289330 294890 289510 294978
rect 289764 294890 289944 294978
rect 290052 294890 290232 294978
rect 290340 294890 290520 294978
rect 290628 294890 290808 294978
rect 290916 294890 291096 294978
rect 291204 294890 291384 294978
rect 291492 294890 291672 294978
rect 291780 294890 291960 294978
rect 292214 294890 292394 294978
rect 292502 294890 292682 294978
rect 292790 294890 292970 294978
rect 293078 294890 293258 294978
rect 293366 294890 293546 294978
rect 293654 294890 293834 294978
rect 293942 294890 294122 294978
rect 294230 294890 294410 294978
rect 294664 294890 294844 294978
rect 294952 294890 295132 294978
rect 295240 294890 295420 294978
rect 295528 294890 295708 294978
rect 295816 294890 295996 294978
rect 296104 294890 296284 294978
rect 296392 294890 296572 294978
rect 296680 294890 296860 294978
rect 297114 294890 297294 294978
rect 297402 294890 297582 294978
rect 297690 294890 297870 294978
rect 297978 294890 298158 294978
rect 298266 294890 298446 294978
rect 298554 294890 298734 294978
rect 298842 294890 299022 294978
rect 299130 294890 299310 294978
rect 299564 294890 299744 294978
rect 299852 294890 300032 294978
rect 300140 294890 300320 294978
rect 300428 294890 300608 294978
rect 300716 294890 300896 294978
rect 301004 294890 301184 294978
rect 301292 294890 301472 294978
rect 301580 294890 301760 294978
rect 302014 294890 302194 294978
rect 302302 294890 302482 294978
rect 302590 294890 302770 294978
rect 302878 294890 303058 294978
rect 303166 294890 303346 294978
rect 303454 294890 303634 294978
rect 303742 294890 303922 294978
rect 304030 294890 304210 294978
rect 304464 294890 304644 294978
rect 304752 294890 304932 294978
rect 305040 294890 305220 294978
rect 305328 294890 305508 294978
rect 305616 294890 305796 294978
rect 305904 294890 306084 294978
rect 306192 294890 306372 294978
rect 306480 294890 306660 294978
rect 306914 294890 307094 294978
rect 307202 294890 307382 294978
rect 307490 294890 307670 294978
rect 307778 294890 307958 294978
rect 308066 294890 308246 294978
rect 308354 294890 308534 294978
rect 308642 294890 308822 294978
rect 308930 294890 309110 294978
rect 309364 294890 309544 294978
rect 309652 294890 309832 294978
rect 309940 294890 310120 294978
rect 310228 294890 310408 294978
rect 310516 294890 310696 294978
rect 310804 294890 310984 294978
rect 311092 294890 311272 294978
rect 311380 294890 311560 294978
rect 311814 294890 311994 294978
rect 312102 294890 312282 294978
rect 312390 294890 312570 294978
rect 312678 294890 312858 294978
rect 312966 294890 313146 294978
rect 313254 294890 313434 294978
rect 313542 294890 313722 294978
rect 313830 294890 314010 294978
rect 314264 294890 314444 294978
rect 314552 294890 314732 294978
rect 314840 294890 315020 294978
rect 315128 294890 315308 294978
rect 315416 294890 315596 294978
rect 315704 294890 315884 294978
rect 315992 294890 316172 294978
rect 316280 294890 316460 294978
rect 316714 294890 316894 294978
rect 317002 294890 317182 294978
rect 317290 294890 317470 294978
rect 317578 294890 317758 294978
rect 317866 294890 318046 294978
rect 318154 294890 318334 294978
rect 318442 294890 318622 294978
rect 318730 294890 318910 294978
rect 319164 294890 319344 294978
rect 319452 294890 319632 294978
rect 319740 294890 319920 294978
rect 320028 294890 320208 294978
rect 320316 294890 320496 294978
rect 320604 294890 320784 294978
rect 320892 294890 321072 294978
rect 321180 294890 321360 294978
rect 321614 294890 321794 294978
rect 321902 294890 322082 294978
rect 322190 294890 322370 294978
rect 322478 294890 322658 294978
rect 322766 294890 322946 294978
rect 323054 294890 323234 294978
rect 323342 294890 323522 294978
rect 323630 294890 323810 294978
rect 324064 294890 324244 294978
rect 324352 294890 324532 294978
rect 324640 294890 324820 294978
rect 324928 294890 325108 294978
rect 325216 294890 325396 294978
rect 325504 294890 325684 294978
rect 325792 294890 325972 294978
rect 326080 294890 326260 294978
rect 326514 294890 326694 294978
rect 326802 294890 326982 294978
rect 327090 294890 327270 294978
rect 327378 294890 327558 294978
rect 327666 294890 327846 294978
rect 327954 294890 328134 294978
rect 328242 294890 328422 294978
rect 328530 294890 328710 294978
rect 328964 294890 329144 294978
rect 329252 294890 329432 294978
rect 329540 294890 329720 294978
rect 329828 294890 330008 294978
rect 330116 294890 330296 294978
rect 330404 294890 330584 294978
rect 330692 294890 330872 294978
rect 330980 294890 331160 294978
rect 331414 294890 331594 294978
rect 331702 294890 331882 294978
rect 331990 294890 332170 294978
rect 332278 294890 332458 294978
rect 332566 294890 332746 294978
rect 332854 294890 333034 294978
rect 333142 294890 333322 294978
rect 333430 294890 333610 294978
rect 333864 294890 334044 294978
rect 334152 294890 334332 294978
rect 334440 294890 334620 294978
rect 334728 294890 334908 294978
rect 335016 294890 335196 294978
rect 335304 294890 335484 294978
rect 335592 294890 335772 294978
rect 335880 294890 336060 294978
rect 336314 294890 336494 294978
rect 336602 294890 336782 294978
rect 336890 294890 337070 294978
rect 337178 294890 337358 294978
rect 337466 294890 337646 294978
rect 337754 294890 337934 294978
rect 338042 294890 338222 294978
rect 338330 294890 338510 294978
rect 338764 294890 338944 294978
rect 339052 294890 339232 294978
rect 339340 294890 339520 294978
rect 339628 294890 339808 294978
rect 339916 294890 340096 294978
rect 340204 294890 340384 294978
rect 340492 294890 340672 294978
rect 340780 294890 340960 294978
rect 341214 294890 341394 294978
rect 341502 294890 341682 294978
rect 341790 294890 341970 294978
rect 342078 294890 342258 294978
rect 342366 294890 342546 294978
rect 342654 294890 342834 294978
rect 342942 294890 343122 294978
rect 343230 294890 343410 294978
rect 343664 294890 343844 294978
rect 343952 294890 344132 294978
rect 344240 294890 344420 294978
rect 344528 294890 344708 294978
rect 344816 294890 344996 294978
rect 345104 294890 345284 294978
rect 345392 294890 345572 294978
rect 345680 294890 345860 294978
rect 346114 294890 346294 294978
rect 346402 294890 346582 294978
rect 346690 294890 346870 294978
rect 346978 294890 347158 294978
rect 347266 294890 347446 294978
rect 347554 294890 347734 294978
rect 347842 294890 348022 294978
rect 348130 294890 348310 294978
rect 348564 294890 348744 294978
rect 348852 294890 349032 294978
rect 349140 294890 349320 294978
rect 349428 294890 349608 294978
rect 349716 294890 349896 294978
rect 350004 294890 350184 294978
rect 350292 294890 350472 294978
rect 350580 294890 350760 294978
rect 351014 294890 351194 294978
rect 351302 294890 351482 294978
rect 351590 294890 351770 294978
rect 351878 294890 352058 294978
rect 352166 294890 352346 294978
rect 352454 294890 352634 294978
rect 352742 294890 352922 294978
rect 353030 294890 353210 294978
rect 353464 294890 353644 294978
rect 353752 294890 353932 294978
rect 354040 294890 354220 294978
rect 354328 294890 354508 294978
rect 354616 294890 354796 294978
rect 354904 294890 355084 294978
rect 355192 294890 355372 294978
rect 355480 294890 355660 294978
rect 355914 294890 356094 294978
rect 356202 294890 356382 294978
rect 356490 294890 356670 294978
rect 356778 294890 356958 294978
rect 357066 294890 357246 294978
rect 357354 294890 357534 294978
rect 357642 294890 357822 294978
rect 357930 294890 358110 294978
rect 358364 294890 358544 294978
rect 358652 294890 358832 294978
rect 358940 294890 359120 294978
rect 359228 294890 359408 294978
rect 359516 294890 359696 294978
rect 359804 294890 359984 294978
rect 360092 294890 360272 294978
rect 360380 294890 360560 294978
rect 360814 294890 360994 294978
rect 361102 294890 361282 294978
rect 361390 294890 361570 294978
rect 361678 294890 361858 294978
rect 361966 294890 362146 294978
rect 362254 294890 362434 294978
rect 362542 294890 362722 294978
rect 362830 294890 363010 294978
rect 363264 294890 363444 294978
rect 363552 294890 363732 294978
rect 363840 294890 364020 294978
rect 364128 294890 364308 294978
rect 364416 294890 364596 294978
rect 364704 294890 364884 294978
rect 364992 294890 365172 294978
rect 365280 294890 365460 294978
rect 365714 294890 365894 294978
rect 366002 294890 366182 294978
rect 366290 294890 366470 294978
rect 366578 294890 366758 294978
rect 366866 294890 367046 294978
rect 367154 294890 367334 294978
rect 367442 294890 367622 294978
rect 367730 294890 367910 294978
rect 243214 294674 243394 294762
rect 243502 294674 243682 294762
rect 243790 294674 243970 294762
rect 244078 294674 244258 294762
rect 244366 294674 244546 294762
rect 244654 294674 244834 294762
rect 244942 294674 245122 294762
rect 245230 294674 245410 294762
rect 245664 294674 245844 294762
rect 245952 294674 246132 294762
rect 246240 294674 246420 294762
rect 246528 294674 246708 294762
rect 246816 294674 246996 294762
rect 247104 294674 247284 294762
rect 247392 294674 247572 294762
rect 247680 294674 247860 294762
rect 248114 294674 248294 294762
rect 248402 294674 248582 294762
rect 248690 294674 248870 294762
rect 248978 294674 249158 294762
rect 249266 294674 249446 294762
rect 249554 294674 249734 294762
rect 249842 294674 250022 294762
rect 250130 294674 250310 294762
rect 250564 294674 250744 294762
rect 250852 294674 251032 294762
rect 251140 294674 251320 294762
rect 251428 294674 251608 294762
rect 251716 294674 251896 294762
rect 252004 294674 252184 294762
rect 252292 294674 252472 294762
rect 252580 294674 252760 294762
rect 253014 294674 253194 294762
rect 253302 294674 253482 294762
rect 253590 294674 253770 294762
rect 253878 294674 254058 294762
rect 254166 294674 254346 294762
rect 254454 294674 254634 294762
rect 254742 294674 254922 294762
rect 255030 294674 255210 294762
rect 255464 294674 255644 294762
rect 255752 294674 255932 294762
rect 256040 294674 256220 294762
rect 256328 294674 256508 294762
rect 256616 294674 256796 294762
rect 256904 294674 257084 294762
rect 257192 294674 257372 294762
rect 257480 294674 257660 294762
rect 257914 294674 258094 294762
rect 258202 294674 258382 294762
rect 258490 294674 258670 294762
rect 258778 294674 258958 294762
rect 259066 294674 259246 294762
rect 259354 294674 259534 294762
rect 259642 294674 259822 294762
rect 259930 294674 260110 294762
rect 260364 294674 260544 294762
rect 260652 294674 260832 294762
rect 260940 294674 261120 294762
rect 261228 294674 261408 294762
rect 261516 294674 261696 294762
rect 261804 294674 261984 294762
rect 262092 294674 262272 294762
rect 262380 294674 262560 294762
rect 262814 294674 262994 294762
rect 263102 294674 263282 294762
rect 263390 294674 263570 294762
rect 263678 294674 263858 294762
rect 263966 294674 264146 294762
rect 264254 294674 264434 294762
rect 264542 294674 264722 294762
rect 264830 294674 265010 294762
rect 265264 294674 265444 294762
rect 265552 294674 265732 294762
rect 265840 294674 266020 294762
rect 266128 294674 266308 294762
rect 266416 294674 266596 294762
rect 266704 294674 266884 294762
rect 266992 294674 267172 294762
rect 267280 294674 267460 294762
rect 267714 294674 267894 294762
rect 268002 294674 268182 294762
rect 268290 294674 268470 294762
rect 268578 294674 268758 294762
rect 268866 294674 269046 294762
rect 269154 294674 269334 294762
rect 269442 294674 269622 294762
rect 269730 294674 269910 294762
rect 270164 294674 270344 294762
rect 270452 294674 270632 294762
rect 270740 294674 270920 294762
rect 271028 294674 271208 294762
rect 271316 294674 271496 294762
rect 271604 294674 271784 294762
rect 271892 294674 272072 294762
rect 272180 294674 272360 294762
rect 272614 294674 272794 294762
rect 272902 294674 273082 294762
rect 273190 294674 273370 294762
rect 273478 294674 273658 294762
rect 273766 294674 273946 294762
rect 274054 294674 274234 294762
rect 274342 294674 274522 294762
rect 274630 294674 274810 294762
rect 275064 294674 275244 294762
rect 275352 294674 275532 294762
rect 275640 294674 275820 294762
rect 275928 294674 276108 294762
rect 276216 294674 276396 294762
rect 276504 294674 276684 294762
rect 276792 294674 276972 294762
rect 277080 294674 277260 294762
rect 277514 294674 277694 294762
rect 277802 294674 277982 294762
rect 278090 294674 278270 294762
rect 278378 294674 278558 294762
rect 278666 294674 278846 294762
rect 278954 294674 279134 294762
rect 279242 294674 279422 294762
rect 279530 294674 279710 294762
rect 279964 294674 280144 294762
rect 280252 294674 280432 294762
rect 280540 294674 280720 294762
rect 280828 294674 281008 294762
rect 281116 294674 281296 294762
rect 281404 294674 281584 294762
rect 281692 294674 281872 294762
rect 281980 294674 282160 294762
rect 282414 294674 282594 294762
rect 282702 294674 282882 294762
rect 282990 294674 283170 294762
rect 283278 294674 283458 294762
rect 283566 294674 283746 294762
rect 283854 294674 284034 294762
rect 284142 294674 284322 294762
rect 284430 294674 284610 294762
rect 284864 294674 285044 294762
rect 285152 294674 285332 294762
rect 285440 294674 285620 294762
rect 285728 294674 285908 294762
rect 286016 294674 286196 294762
rect 286304 294674 286484 294762
rect 286592 294674 286772 294762
rect 286880 294674 287060 294762
rect 287314 294674 287494 294762
rect 287602 294674 287782 294762
rect 287890 294674 288070 294762
rect 288178 294674 288358 294762
rect 288466 294674 288646 294762
rect 288754 294674 288934 294762
rect 289042 294674 289222 294762
rect 289330 294674 289510 294762
rect 289764 294674 289944 294762
rect 290052 294674 290232 294762
rect 290340 294674 290520 294762
rect 290628 294674 290808 294762
rect 290916 294674 291096 294762
rect 291204 294674 291384 294762
rect 291492 294674 291672 294762
rect 291780 294674 291960 294762
rect 292214 294674 292394 294762
rect 292502 294674 292682 294762
rect 292790 294674 292970 294762
rect 293078 294674 293258 294762
rect 293366 294674 293546 294762
rect 293654 294674 293834 294762
rect 293942 294674 294122 294762
rect 294230 294674 294410 294762
rect 294664 294674 294844 294762
rect 294952 294674 295132 294762
rect 295240 294674 295420 294762
rect 295528 294674 295708 294762
rect 295816 294674 295996 294762
rect 296104 294674 296284 294762
rect 296392 294674 296572 294762
rect 296680 294674 296860 294762
rect 297114 294674 297294 294762
rect 297402 294674 297582 294762
rect 297690 294674 297870 294762
rect 297978 294674 298158 294762
rect 298266 294674 298446 294762
rect 298554 294674 298734 294762
rect 298842 294674 299022 294762
rect 299130 294674 299310 294762
rect 299564 294674 299744 294762
rect 299852 294674 300032 294762
rect 300140 294674 300320 294762
rect 300428 294674 300608 294762
rect 300716 294674 300896 294762
rect 301004 294674 301184 294762
rect 301292 294674 301472 294762
rect 301580 294674 301760 294762
rect 302014 294674 302194 294762
rect 302302 294674 302482 294762
rect 302590 294674 302770 294762
rect 302878 294674 303058 294762
rect 303166 294674 303346 294762
rect 303454 294674 303634 294762
rect 303742 294674 303922 294762
rect 304030 294674 304210 294762
rect 304464 294674 304644 294762
rect 304752 294674 304932 294762
rect 305040 294674 305220 294762
rect 305328 294674 305508 294762
rect 305616 294674 305796 294762
rect 305904 294674 306084 294762
rect 306192 294674 306372 294762
rect 306480 294674 306660 294762
rect 306914 294674 307094 294762
rect 307202 294674 307382 294762
rect 307490 294674 307670 294762
rect 307778 294674 307958 294762
rect 308066 294674 308246 294762
rect 308354 294674 308534 294762
rect 308642 294674 308822 294762
rect 308930 294674 309110 294762
rect 309364 294674 309544 294762
rect 309652 294674 309832 294762
rect 309940 294674 310120 294762
rect 310228 294674 310408 294762
rect 310516 294674 310696 294762
rect 310804 294674 310984 294762
rect 311092 294674 311272 294762
rect 311380 294674 311560 294762
rect 311814 294674 311994 294762
rect 312102 294674 312282 294762
rect 312390 294674 312570 294762
rect 312678 294674 312858 294762
rect 312966 294674 313146 294762
rect 313254 294674 313434 294762
rect 313542 294674 313722 294762
rect 313830 294674 314010 294762
rect 314264 294674 314444 294762
rect 314552 294674 314732 294762
rect 314840 294674 315020 294762
rect 315128 294674 315308 294762
rect 315416 294674 315596 294762
rect 315704 294674 315884 294762
rect 315992 294674 316172 294762
rect 316280 294674 316460 294762
rect 316714 294674 316894 294762
rect 317002 294674 317182 294762
rect 317290 294674 317470 294762
rect 317578 294674 317758 294762
rect 317866 294674 318046 294762
rect 318154 294674 318334 294762
rect 318442 294674 318622 294762
rect 318730 294674 318910 294762
rect 319164 294674 319344 294762
rect 319452 294674 319632 294762
rect 319740 294674 319920 294762
rect 320028 294674 320208 294762
rect 320316 294674 320496 294762
rect 320604 294674 320784 294762
rect 320892 294674 321072 294762
rect 321180 294674 321360 294762
rect 321614 294674 321794 294762
rect 321902 294674 322082 294762
rect 322190 294674 322370 294762
rect 322478 294674 322658 294762
rect 322766 294674 322946 294762
rect 323054 294674 323234 294762
rect 323342 294674 323522 294762
rect 323630 294674 323810 294762
rect 324064 294674 324244 294762
rect 324352 294674 324532 294762
rect 324640 294674 324820 294762
rect 324928 294674 325108 294762
rect 325216 294674 325396 294762
rect 325504 294674 325684 294762
rect 325792 294674 325972 294762
rect 326080 294674 326260 294762
rect 326514 294674 326694 294762
rect 326802 294674 326982 294762
rect 327090 294674 327270 294762
rect 327378 294674 327558 294762
rect 327666 294674 327846 294762
rect 327954 294674 328134 294762
rect 328242 294674 328422 294762
rect 328530 294674 328710 294762
rect 328964 294674 329144 294762
rect 329252 294674 329432 294762
rect 329540 294674 329720 294762
rect 329828 294674 330008 294762
rect 330116 294674 330296 294762
rect 330404 294674 330584 294762
rect 330692 294674 330872 294762
rect 330980 294674 331160 294762
rect 331414 294674 331594 294762
rect 331702 294674 331882 294762
rect 331990 294674 332170 294762
rect 332278 294674 332458 294762
rect 332566 294674 332746 294762
rect 332854 294674 333034 294762
rect 333142 294674 333322 294762
rect 333430 294674 333610 294762
rect 333864 294674 334044 294762
rect 334152 294674 334332 294762
rect 334440 294674 334620 294762
rect 334728 294674 334908 294762
rect 335016 294674 335196 294762
rect 335304 294674 335484 294762
rect 335592 294674 335772 294762
rect 335880 294674 336060 294762
rect 336314 294674 336494 294762
rect 336602 294674 336782 294762
rect 336890 294674 337070 294762
rect 337178 294674 337358 294762
rect 337466 294674 337646 294762
rect 337754 294674 337934 294762
rect 338042 294674 338222 294762
rect 338330 294674 338510 294762
rect 338764 294674 338944 294762
rect 339052 294674 339232 294762
rect 339340 294674 339520 294762
rect 339628 294674 339808 294762
rect 339916 294674 340096 294762
rect 340204 294674 340384 294762
rect 340492 294674 340672 294762
rect 340780 294674 340960 294762
rect 341214 294674 341394 294762
rect 341502 294674 341682 294762
rect 341790 294674 341970 294762
rect 342078 294674 342258 294762
rect 342366 294674 342546 294762
rect 342654 294674 342834 294762
rect 342942 294674 343122 294762
rect 343230 294674 343410 294762
rect 343664 294674 343844 294762
rect 343952 294674 344132 294762
rect 344240 294674 344420 294762
rect 344528 294674 344708 294762
rect 344816 294674 344996 294762
rect 345104 294674 345284 294762
rect 345392 294674 345572 294762
rect 345680 294674 345860 294762
rect 346114 294674 346294 294762
rect 346402 294674 346582 294762
rect 346690 294674 346870 294762
rect 346978 294674 347158 294762
rect 347266 294674 347446 294762
rect 347554 294674 347734 294762
rect 347842 294674 348022 294762
rect 348130 294674 348310 294762
rect 348564 294674 348744 294762
rect 348852 294674 349032 294762
rect 349140 294674 349320 294762
rect 349428 294674 349608 294762
rect 349716 294674 349896 294762
rect 350004 294674 350184 294762
rect 350292 294674 350472 294762
rect 350580 294674 350760 294762
rect 351014 294674 351194 294762
rect 351302 294674 351482 294762
rect 351590 294674 351770 294762
rect 351878 294674 352058 294762
rect 352166 294674 352346 294762
rect 352454 294674 352634 294762
rect 352742 294674 352922 294762
rect 353030 294674 353210 294762
rect 353464 294674 353644 294762
rect 353752 294674 353932 294762
rect 354040 294674 354220 294762
rect 354328 294674 354508 294762
rect 354616 294674 354796 294762
rect 354904 294674 355084 294762
rect 355192 294674 355372 294762
rect 355480 294674 355660 294762
rect 355914 294674 356094 294762
rect 356202 294674 356382 294762
rect 356490 294674 356670 294762
rect 356778 294674 356958 294762
rect 357066 294674 357246 294762
rect 357354 294674 357534 294762
rect 357642 294674 357822 294762
rect 357930 294674 358110 294762
rect 358364 294674 358544 294762
rect 358652 294674 358832 294762
rect 358940 294674 359120 294762
rect 359228 294674 359408 294762
rect 359516 294674 359696 294762
rect 359804 294674 359984 294762
rect 360092 294674 360272 294762
rect 360380 294674 360560 294762
rect 360814 294674 360994 294762
rect 361102 294674 361282 294762
rect 361390 294674 361570 294762
rect 361678 294674 361858 294762
rect 361966 294674 362146 294762
rect 362254 294674 362434 294762
rect 362542 294674 362722 294762
rect 362830 294674 363010 294762
rect 363264 294674 363444 294762
rect 363552 294674 363732 294762
rect 363840 294674 364020 294762
rect 364128 294674 364308 294762
rect 364416 294674 364596 294762
rect 364704 294674 364884 294762
rect 364992 294674 365172 294762
rect 365280 294674 365460 294762
rect 365714 294674 365894 294762
rect 366002 294674 366182 294762
rect 366290 294674 366470 294762
rect 366578 294674 366758 294762
rect 366866 294674 367046 294762
rect 367154 294674 367334 294762
rect 367442 294674 367622 294762
rect 367730 294674 367910 294762
rect 243214 294198 243394 294286
rect 243502 294198 243682 294286
rect 243790 294198 243970 294286
rect 244078 294198 244258 294286
rect 244366 294198 244546 294286
rect 244654 294198 244834 294286
rect 244942 294198 245122 294286
rect 245230 294198 245410 294286
rect 245664 294198 245844 294286
rect 245952 294198 246132 294286
rect 246240 294198 246420 294286
rect 246528 294198 246708 294286
rect 246816 294198 246996 294286
rect 247104 294198 247284 294286
rect 247392 294198 247572 294286
rect 247680 294198 247860 294286
rect 248114 294198 248294 294286
rect 248402 294198 248582 294286
rect 248690 294198 248870 294286
rect 248978 294198 249158 294286
rect 249266 294198 249446 294286
rect 249554 294198 249734 294286
rect 249842 294198 250022 294286
rect 250130 294198 250310 294286
rect 250564 294198 250744 294286
rect 250852 294198 251032 294286
rect 251140 294198 251320 294286
rect 251428 294198 251608 294286
rect 251716 294198 251896 294286
rect 252004 294198 252184 294286
rect 252292 294198 252472 294286
rect 252580 294198 252760 294286
rect 253014 294198 253194 294286
rect 253302 294198 253482 294286
rect 253590 294198 253770 294286
rect 253878 294198 254058 294286
rect 254166 294198 254346 294286
rect 254454 294198 254634 294286
rect 254742 294198 254922 294286
rect 255030 294198 255210 294286
rect 255464 294198 255644 294286
rect 255752 294198 255932 294286
rect 256040 294198 256220 294286
rect 256328 294198 256508 294286
rect 256616 294198 256796 294286
rect 256904 294198 257084 294286
rect 257192 294198 257372 294286
rect 257480 294198 257660 294286
rect 257914 294198 258094 294286
rect 258202 294198 258382 294286
rect 258490 294198 258670 294286
rect 258778 294198 258958 294286
rect 259066 294198 259246 294286
rect 259354 294198 259534 294286
rect 259642 294198 259822 294286
rect 259930 294198 260110 294286
rect 260364 294198 260544 294286
rect 260652 294198 260832 294286
rect 260940 294198 261120 294286
rect 261228 294198 261408 294286
rect 261516 294198 261696 294286
rect 261804 294198 261984 294286
rect 262092 294198 262272 294286
rect 262380 294198 262560 294286
rect 262814 294198 262994 294286
rect 263102 294198 263282 294286
rect 263390 294198 263570 294286
rect 263678 294198 263858 294286
rect 263966 294198 264146 294286
rect 264254 294198 264434 294286
rect 264542 294198 264722 294286
rect 264830 294198 265010 294286
rect 265264 294198 265444 294286
rect 265552 294198 265732 294286
rect 265840 294198 266020 294286
rect 266128 294198 266308 294286
rect 266416 294198 266596 294286
rect 266704 294198 266884 294286
rect 266992 294198 267172 294286
rect 267280 294198 267460 294286
rect 267714 294198 267894 294286
rect 268002 294198 268182 294286
rect 268290 294198 268470 294286
rect 268578 294198 268758 294286
rect 268866 294198 269046 294286
rect 269154 294198 269334 294286
rect 269442 294198 269622 294286
rect 269730 294198 269910 294286
rect 270164 294198 270344 294286
rect 270452 294198 270632 294286
rect 270740 294198 270920 294286
rect 271028 294198 271208 294286
rect 271316 294198 271496 294286
rect 271604 294198 271784 294286
rect 271892 294198 272072 294286
rect 272180 294198 272360 294286
rect 272614 294198 272794 294286
rect 272902 294198 273082 294286
rect 273190 294198 273370 294286
rect 273478 294198 273658 294286
rect 273766 294198 273946 294286
rect 274054 294198 274234 294286
rect 274342 294198 274522 294286
rect 274630 294198 274810 294286
rect 275064 294198 275244 294286
rect 275352 294198 275532 294286
rect 275640 294198 275820 294286
rect 275928 294198 276108 294286
rect 276216 294198 276396 294286
rect 276504 294198 276684 294286
rect 276792 294198 276972 294286
rect 277080 294198 277260 294286
rect 277514 294198 277694 294286
rect 277802 294198 277982 294286
rect 278090 294198 278270 294286
rect 278378 294198 278558 294286
rect 278666 294198 278846 294286
rect 278954 294198 279134 294286
rect 279242 294198 279422 294286
rect 279530 294198 279710 294286
rect 279964 294198 280144 294286
rect 280252 294198 280432 294286
rect 280540 294198 280720 294286
rect 280828 294198 281008 294286
rect 281116 294198 281296 294286
rect 281404 294198 281584 294286
rect 281692 294198 281872 294286
rect 281980 294198 282160 294286
rect 282414 294198 282594 294286
rect 282702 294198 282882 294286
rect 282990 294198 283170 294286
rect 283278 294198 283458 294286
rect 283566 294198 283746 294286
rect 283854 294198 284034 294286
rect 284142 294198 284322 294286
rect 284430 294198 284610 294286
rect 284864 294198 285044 294286
rect 285152 294198 285332 294286
rect 285440 294198 285620 294286
rect 285728 294198 285908 294286
rect 286016 294198 286196 294286
rect 286304 294198 286484 294286
rect 286592 294198 286772 294286
rect 286880 294198 287060 294286
rect 287314 294198 287494 294286
rect 287602 294198 287782 294286
rect 287890 294198 288070 294286
rect 288178 294198 288358 294286
rect 288466 294198 288646 294286
rect 288754 294198 288934 294286
rect 289042 294198 289222 294286
rect 289330 294198 289510 294286
rect 289764 294198 289944 294286
rect 290052 294198 290232 294286
rect 290340 294198 290520 294286
rect 290628 294198 290808 294286
rect 290916 294198 291096 294286
rect 291204 294198 291384 294286
rect 291492 294198 291672 294286
rect 291780 294198 291960 294286
rect 292214 294198 292394 294286
rect 292502 294198 292682 294286
rect 292790 294198 292970 294286
rect 293078 294198 293258 294286
rect 293366 294198 293546 294286
rect 293654 294198 293834 294286
rect 293942 294198 294122 294286
rect 294230 294198 294410 294286
rect 294664 294198 294844 294286
rect 294952 294198 295132 294286
rect 295240 294198 295420 294286
rect 295528 294198 295708 294286
rect 295816 294198 295996 294286
rect 296104 294198 296284 294286
rect 296392 294198 296572 294286
rect 296680 294198 296860 294286
rect 297114 294198 297294 294286
rect 297402 294198 297582 294286
rect 297690 294198 297870 294286
rect 297978 294198 298158 294286
rect 298266 294198 298446 294286
rect 298554 294198 298734 294286
rect 298842 294198 299022 294286
rect 299130 294198 299310 294286
rect 299564 294198 299744 294286
rect 299852 294198 300032 294286
rect 300140 294198 300320 294286
rect 300428 294198 300608 294286
rect 300716 294198 300896 294286
rect 301004 294198 301184 294286
rect 301292 294198 301472 294286
rect 301580 294198 301760 294286
rect 302014 294198 302194 294286
rect 302302 294198 302482 294286
rect 302590 294198 302770 294286
rect 302878 294198 303058 294286
rect 303166 294198 303346 294286
rect 303454 294198 303634 294286
rect 303742 294198 303922 294286
rect 304030 294198 304210 294286
rect 304464 294198 304644 294286
rect 304752 294198 304932 294286
rect 305040 294198 305220 294286
rect 305328 294198 305508 294286
rect 305616 294198 305796 294286
rect 305904 294198 306084 294286
rect 306192 294198 306372 294286
rect 306480 294198 306660 294286
rect 306914 294198 307094 294286
rect 307202 294198 307382 294286
rect 307490 294198 307670 294286
rect 307778 294198 307958 294286
rect 308066 294198 308246 294286
rect 308354 294198 308534 294286
rect 308642 294198 308822 294286
rect 308930 294198 309110 294286
rect 309364 294198 309544 294286
rect 309652 294198 309832 294286
rect 309940 294198 310120 294286
rect 310228 294198 310408 294286
rect 310516 294198 310696 294286
rect 310804 294198 310984 294286
rect 311092 294198 311272 294286
rect 311380 294198 311560 294286
rect 311814 294198 311994 294286
rect 312102 294198 312282 294286
rect 312390 294198 312570 294286
rect 312678 294198 312858 294286
rect 312966 294198 313146 294286
rect 313254 294198 313434 294286
rect 313542 294198 313722 294286
rect 313830 294198 314010 294286
rect 314264 294198 314444 294286
rect 314552 294198 314732 294286
rect 314840 294198 315020 294286
rect 315128 294198 315308 294286
rect 315416 294198 315596 294286
rect 315704 294198 315884 294286
rect 315992 294198 316172 294286
rect 316280 294198 316460 294286
rect 316714 294198 316894 294286
rect 317002 294198 317182 294286
rect 317290 294198 317470 294286
rect 317578 294198 317758 294286
rect 317866 294198 318046 294286
rect 318154 294198 318334 294286
rect 318442 294198 318622 294286
rect 318730 294198 318910 294286
rect 319164 294198 319344 294286
rect 319452 294198 319632 294286
rect 319740 294198 319920 294286
rect 320028 294198 320208 294286
rect 320316 294198 320496 294286
rect 320604 294198 320784 294286
rect 320892 294198 321072 294286
rect 321180 294198 321360 294286
rect 321614 294198 321794 294286
rect 321902 294198 322082 294286
rect 322190 294198 322370 294286
rect 322478 294198 322658 294286
rect 322766 294198 322946 294286
rect 323054 294198 323234 294286
rect 323342 294198 323522 294286
rect 323630 294198 323810 294286
rect 324064 294198 324244 294286
rect 324352 294198 324532 294286
rect 324640 294198 324820 294286
rect 324928 294198 325108 294286
rect 325216 294198 325396 294286
rect 325504 294198 325684 294286
rect 325792 294198 325972 294286
rect 326080 294198 326260 294286
rect 326514 294198 326694 294286
rect 326802 294198 326982 294286
rect 327090 294198 327270 294286
rect 327378 294198 327558 294286
rect 327666 294198 327846 294286
rect 327954 294198 328134 294286
rect 328242 294198 328422 294286
rect 328530 294198 328710 294286
rect 328964 294198 329144 294286
rect 329252 294198 329432 294286
rect 329540 294198 329720 294286
rect 329828 294198 330008 294286
rect 330116 294198 330296 294286
rect 330404 294198 330584 294286
rect 330692 294198 330872 294286
rect 330980 294198 331160 294286
rect 331414 294198 331594 294286
rect 331702 294198 331882 294286
rect 331990 294198 332170 294286
rect 332278 294198 332458 294286
rect 332566 294198 332746 294286
rect 332854 294198 333034 294286
rect 333142 294198 333322 294286
rect 333430 294198 333610 294286
rect 333864 294198 334044 294286
rect 334152 294198 334332 294286
rect 334440 294198 334620 294286
rect 334728 294198 334908 294286
rect 335016 294198 335196 294286
rect 335304 294198 335484 294286
rect 335592 294198 335772 294286
rect 335880 294198 336060 294286
rect 336314 294198 336494 294286
rect 336602 294198 336782 294286
rect 336890 294198 337070 294286
rect 337178 294198 337358 294286
rect 337466 294198 337646 294286
rect 337754 294198 337934 294286
rect 338042 294198 338222 294286
rect 338330 294198 338510 294286
rect 338764 294198 338944 294286
rect 339052 294198 339232 294286
rect 339340 294198 339520 294286
rect 339628 294198 339808 294286
rect 339916 294198 340096 294286
rect 340204 294198 340384 294286
rect 340492 294198 340672 294286
rect 340780 294198 340960 294286
rect 341214 294198 341394 294286
rect 341502 294198 341682 294286
rect 341790 294198 341970 294286
rect 342078 294198 342258 294286
rect 342366 294198 342546 294286
rect 342654 294198 342834 294286
rect 342942 294198 343122 294286
rect 343230 294198 343410 294286
rect 343664 294198 343844 294286
rect 343952 294198 344132 294286
rect 344240 294198 344420 294286
rect 344528 294198 344708 294286
rect 344816 294198 344996 294286
rect 345104 294198 345284 294286
rect 345392 294198 345572 294286
rect 345680 294198 345860 294286
rect 346114 294198 346294 294286
rect 346402 294198 346582 294286
rect 346690 294198 346870 294286
rect 346978 294198 347158 294286
rect 347266 294198 347446 294286
rect 347554 294198 347734 294286
rect 347842 294198 348022 294286
rect 348130 294198 348310 294286
rect 348564 294198 348744 294286
rect 348852 294198 349032 294286
rect 349140 294198 349320 294286
rect 349428 294198 349608 294286
rect 349716 294198 349896 294286
rect 350004 294198 350184 294286
rect 350292 294198 350472 294286
rect 350580 294198 350760 294286
rect 351014 294198 351194 294286
rect 351302 294198 351482 294286
rect 351590 294198 351770 294286
rect 351878 294198 352058 294286
rect 352166 294198 352346 294286
rect 352454 294198 352634 294286
rect 352742 294198 352922 294286
rect 353030 294198 353210 294286
rect 353464 294198 353644 294286
rect 353752 294198 353932 294286
rect 354040 294198 354220 294286
rect 354328 294198 354508 294286
rect 354616 294198 354796 294286
rect 354904 294198 355084 294286
rect 355192 294198 355372 294286
rect 355480 294198 355660 294286
rect 355914 294198 356094 294286
rect 356202 294198 356382 294286
rect 356490 294198 356670 294286
rect 356778 294198 356958 294286
rect 357066 294198 357246 294286
rect 357354 294198 357534 294286
rect 357642 294198 357822 294286
rect 357930 294198 358110 294286
rect 358364 294198 358544 294286
rect 358652 294198 358832 294286
rect 358940 294198 359120 294286
rect 359228 294198 359408 294286
rect 359516 294198 359696 294286
rect 359804 294198 359984 294286
rect 360092 294198 360272 294286
rect 360380 294198 360560 294286
rect 360814 294198 360994 294286
rect 361102 294198 361282 294286
rect 361390 294198 361570 294286
rect 361678 294198 361858 294286
rect 361966 294198 362146 294286
rect 362254 294198 362434 294286
rect 362542 294198 362722 294286
rect 362830 294198 363010 294286
rect 363264 294198 363444 294286
rect 363552 294198 363732 294286
rect 363840 294198 364020 294286
rect 364128 294198 364308 294286
rect 364416 294198 364596 294286
rect 364704 294198 364884 294286
rect 364992 294198 365172 294286
rect 365280 294198 365460 294286
rect 365714 294198 365894 294286
rect 366002 294198 366182 294286
rect 366290 294198 366470 294286
rect 366578 294198 366758 294286
rect 366866 294198 367046 294286
rect 367154 294198 367334 294286
rect 367442 294198 367622 294286
rect 367730 294198 367910 294286
rect 243214 293724 243394 293812
rect 243502 293724 243682 293812
rect 243790 293724 243970 293812
rect 244078 293724 244258 293812
rect 244366 293724 244546 293812
rect 244654 293724 244834 293812
rect 244942 293724 245122 293812
rect 245230 293724 245410 293812
rect 245664 293724 245844 293812
rect 245952 293724 246132 293812
rect 246240 293724 246420 293812
rect 246528 293724 246708 293812
rect 246816 293724 246996 293812
rect 247104 293724 247284 293812
rect 247392 293724 247572 293812
rect 247680 293724 247860 293812
rect 248114 293724 248294 293812
rect 248402 293724 248582 293812
rect 248690 293724 248870 293812
rect 248978 293724 249158 293812
rect 249266 293724 249446 293812
rect 249554 293724 249734 293812
rect 249842 293724 250022 293812
rect 250130 293724 250310 293812
rect 250564 293724 250744 293812
rect 250852 293724 251032 293812
rect 251140 293724 251320 293812
rect 251428 293724 251608 293812
rect 251716 293724 251896 293812
rect 252004 293724 252184 293812
rect 252292 293724 252472 293812
rect 252580 293724 252760 293812
rect 253014 293724 253194 293812
rect 253302 293724 253482 293812
rect 253590 293724 253770 293812
rect 253878 293724 254058 293812
rect 254166 293724 254346 293812
rect 254454 293724 254634 293812
rect 254742 293724 254922 293812
rect 255030 293724 255210 293812
rect 255464 293724 255644 293812
rect 255752 293724 255932 293812
rect 256040 293724 256220 293812
rect 256328 293724 256508 293812
rect 256616 293724 256796 293812
rect 256904 293724 257084 293812
rect 257192 293724 257372 293812
rect 257480 293724 257660 293812
rect 257914 293724 258094 293812
rect 258202 293724 258382 293812
rect 258490 293724 258670 293812
rect 258778 293724 258958 293812
rect 259066 293724 259246 293812
rect 259354 293724 259534 293812
rect 259642 293724 259822 293812
rect 259930 293724 260110 293812
rect 260364 293724 260544 293812
rect 260652 293724 260832 293812
rect 260940 293724 261120 293812
rect 261228 293724 261408 293812
rect 261516 293724 261696 293812
rect 261804 293724 261984 293812
rect 262092 293724 262272 293812
rect 262380 293724 262560 293812
rect 262814 293724 262994 293812
rect 263102 293724 263282 293812
rect 263390 293724 263570 293812
rect 263678 293724 263858 293812
rect 263966 293724 264146 293812
rect 264254 293724 264434 293812
rect 264542 293724 264722 293812
rect 264830 293724 265010 293812
rect 265264 293724 265444 293812
rect 265552 293724 265732 293812
rect 265840 293724 266020 293812
rect 266128 293724 266308 293812
rect 266416 293724 266596 293812
rect 266704 293724 266884 293812
rect 266992 293724 267172 293812
rect 267280 293724 267460 293812
rect 267714 293724 267894 293812
rect 268002 293724 268182 293812
rect 268290 293724 268470 293812
rect 268578 293724 268758 293812
rect 268866 293724 269046 293812
rect 269154 293724 269334 293812
rect 269442 293724 269622 293812
rect 269730 293724 269910 293812
rect 270164 293724 270344 293812
rect 270452 293724 270632 293812
rect 270740 293724 270920 293812
rect 271028 293724 271208 293812
rect 271316 293724 271496 293812
rect 271604 293724 271784 293812
rect 271892 293724 272072 293812
rect 272180 293724 272360 293812
rect 272614 293724 272794 293812
rect 272902 293724 273082 293812
rect 273190 293724 273370 293812
rect 273478 293724 273658 293812
rect 273766 293724 273946 293812
rect 274054 293724 274234 293812
rect 274342 293724 274522 293812
rect 274630 293724 274810 293812
rect 275064 293724 275244 293812
rect 275352 293724 275532 293812
rect 275640 293724 275820 293812
rect 275928 293724 276108 293812
rect 276216 293724 276396 293812
rect 276504 293724 276684 293812
rect 276792 293724 276972 293812
rect 277080 293724 277260 293812
rect 277514 293724 277694 293812
rect 277802 293724 277982 293812
rect 278090 293724 278270 293812
rect 278378 293724 278558 293812
rect 278666 293724 278846 293812
rect 278954 293724 279134 293812
rect 279242 293724 279422 293812
rect 279530 293724 279710 293812
rect 279964 293724 280144 293812
rect 280252 293724 280432 293812
rect 280540 293724 280720 293812
rect 280828 293724 281008 293812
rect 281116 293724 281296 293812
rect 281404 293724 281584 293812
rect 281692 293724 281872 293812
rect 281980 293724 282160 293812
rect 282414 293724 282594 293812
rect 282702 293724 282882 293812
rect 282990 293724 283170 293812
rect 283278 293724 283458 293812
rect 283566 293724 283746 293812
rect 283854 293724 284034 293812
rect 284142 293724 284322 293812
rect 284430 293724 284610 293812
rect 284864 293724 285044 293812
rect 285152 293724 285332 293812
rect 285440 293724 285620 293812
rect 285728 293724 285908 293812
rect 286016 293724 286196 293812
rect 286304 293724 286484 293812
rect 286592 293724 286772 293812
rect 286880 293724 287060 293812
rect 287314 293724 287494 293812
rect 287602 293724 287782 293812
rect 287890 293724 288070 293812
rect 288178 293724 288358 293812
rect 288466 293724 288646 293812
rect 288754 293724 288934 293812
rect 289042 293724 289222 293812
rect 289330 293724 289510 293812
rect 289764 293724 289944 293812
rect 290052 293724 290232 293812
rect 290340 293724 290520 293812
rect 290628 293724 290808 293812
rect 290916 293724 291096 293812
rect 291204 293724 291384 293812
rect 291492 293724 291672 293812
rect 291780 293724 291960 293812
rect 292214 293724 292394 293812
rect 292502 293724 292682 293812
rect 292790 293724 292970 293812
rect 293078 293724 293258 293812
rect 293366 293724 293546 293812
rect 293654 293724 293834 293812
rect 293942 293724 294122 293812
rect 294230 293724 294410 293812
rect 294664 293724 294844 293812
rect 294952 293724 295132 293812
rect 295240 293724 295420 293812
rect 295528 293724 295708 293812
rect 295816 293724 295996 293812
rect 296104 293724 296284 293812
rect 296392 293724 296572 293812
rect 296680 293724 296860 293812
rect 297114 293724 297294 293812
rect 297402 293724 297582 293812
rect 297690 293724 297870 293812
rect 297978 293724 298158 293812
rect 298266 293724 298446 293812
rect 298554 293724 298734 293812
rect 298842 293724 299022 293812
rect 299130 293724 299310 293812
rect 299564 293724 299744 293812
rect 299852 293724 300032 293812
rect 300140 293724 300320 293812
rect 300428 293724 300608 293812
rect 300716 293724 300896 293812
rect 301004 293724 301184 293812
rect 301292 293724 301472 293812
rect 301580 293724 301760 293812
rect 302014 293724 302194 293812
rect 302302 293724 302482 293812
rect 302590 293724 302770 293812
rect 302878 293724 303058 293812
rect 303166 293724 303346 293812
rect 303454 293724 303634 293812
rect 303742 293724 303922 293812
rect 304030 293724 304210 293812
rect 304464 293724 304644 293812
rect 304752 293724 304932 293812
rect 305040 293724 305220 293812
rect 305328 293724 305508 293812
rect 305616 293724 305796 293812
rect 305904 293724 306084 293812
rect 306192 293724 306372 293812
rect 306480 293724 306660 293812
rect 306914 293724 307094 293812
rect 307202 293724 307382 293812
rect 307490 293724 307670 293812
rect 307778 293724 307958 293812
rect 308066 293724 308246 293812
rect 308354 293724 308534 293812
rect 308642 293724 308822 293812
rect 308930 293724 309110 293812
rect 309364 293724 309544 293812
rect 309652 293724 309832 293812
rect 309940 293724 310120 293812
rect 310228 293724 310408 293812
rect 310516 293724 310696 293812
rect 310804 293724 310984 293812
rect 311092 293724 311272 293812
rect 311380 293724 311560 293812
rect 311814 293724 311994 293812
rect 312102 293724 312282 293812
rect 312390 293724 312570 293812
rect 312678 293724 312858 293812
rect 312966 293724 313146 293812
rect 313254 293724 313434 293812
rect 313542 293724 313722 293812
rect 313830 293724 314010 293812
rect 314264 293724 314444 293812
rect 314552 293724 314732 293812
rect 314840 293724 315020 293812
rect 315128 293724 315308 293812
rect 315416 293724 315596 293812
rect 315704 293724 315884 293812
rect 315992 293724 316172 293812
rect 316280 293724 316460 293812
rect 316714 293724 316894 293812
rect 317002 293724 317182 293812
rect 317290 293724 317470 293812
rect 317578 293724 317758 293812
rect 317866 293724 318046 293812
rect 318154 293724 318334 293812
rect 318442 293724 318622 293812
rect 318730 293724 318910 293812
rect 319164 293724 319344 293812
rect 319452 293724 319632 293812
rect 319740 293724 319920 293812
rect 320028 293724 320208 293812
rect 320316 293724 320496 293812
rect 320604 293724 320784 293812
rect 320892 293724 321072 293812
rect 321180 293724 321360 293812
rect 321614 293724 321794 293812
rect 321902 293724 322082 293812
rect 322190 293724 322370 293812
rect 322478 293724 322658 293812
rect 322766 293724 322946 293812
rect 323054 293724 323234 293812
rect 323342 293724 323522 293812
rect 323630 293724 323810 293812
rect 324064 293724 324244 293812
rect 324352 293724 324532 293812
rect 324640 293724 324820 293812
rect 324928 293724 325108 293812
rect 325216 293724 325396 293812
rect 325504 293724 325684 293812
rect 325792 293724 325972 293812
rect 326080 293724 326260 293812
rect 326514 293724 326694 293812
rect 326802 293724 326982 293812
rect 327090 293724 327270 293812
rect 327378 293724 327558 293812
rect 327666 293724 327846 293812
rect 327954 293724 328134 293812
rect 328242 293724 328422 293812
rect 328530 293724 328710 293812
rect 328964 293724 329144 293812
rect 329252 293724 329432 293812
rect 329540 293724 329720 293812
rect 329828 293724 330008 293812
rect 330116 293724 330296 293812
rect 330404 293724 330584 293812
rect 330692 293724 330872 293812
rect 330980 293724 331160 293812
rect 331414 293724 331594 293812
rect 331702 293724 331882 293812
rect 331990 293724 332170 293812
rect 332278 293724 332458 293812
rect 332566 293724 332746 293812
rect 332854 293724 333034 293812
rect 333142 293724 333322 293812
rect 333430 293724 333610 293812
rect 333864 293724 334044 293812
rect 334152 293724 334332 293812
rect 334440 293724 334620 293812
rect 334728 293724 334908 293812
rect 335016 293724 335196 293812
rect 335304 293724 335484 293812
rect 335592 293724 335772 293812
rect 335880 293724 336060 293812
rect 336314 293724 336494 293812
rect 336602 293724 336782 293812
rect 336890 293724 337070 293812
rect 337178 293724 337358 293812
rect 337466 293724 337646 293812
rect 337754 293724 337934 293812
rect 338042 293724 338222 293812
rect 338330 293724 338510 293812
rect 338764 293724 338944 293812
rect 339052 293724 339232 293812
rect 339340 293724 339520 293812
rect 339628 293724 339808 293812
rect 339916 293724 340096 293812
rect 340204 293724 340384 293812
rect 340492 293724 340672 293812
rect 340780 293724 340960 293812
rect 341214 293724 341394 293812
rect 341502 293724 341682 293812
rect 341790 293724 341970 293812
rect 342078 293724 342258 293812
rect 342366 293724 342546 293812
rect 342654 293724 342834 293812
rect 342942 293724 343122 293812
rect 343230 293724 343410 293812
rect 343664 293724 343844 293812
rect 343952 293724 344132 293812
rect 344240 293724 344420 293812
rect 344528 293724 344708 293812
rect 344816 293724 344996 293812
rect 345104 293724 345284 293812
rect 345392 293724 345572 293812
rect 345680 293724 345860 293812
rect 346114 293724 346294 293812
rect 346402 293724 346582 293812
rect 346690 293724 346870 293812
rect 346978 293724 347158 293812
rect 347266 293724 347446 293812
rect 347554 293724 347734 293812
rect 347842 293724 348022 293812
rect 348130 293724 348310 293812
rect 348564 293724 348744 293812
rect 348852 293724 349032 293812
rect 349140 293724 349320 293812
rect 349428 293724 349608 293812
rect 349716 293724 349896 293812
rect 350004 293724 350184 293812
rect 350292 293724 350472 293812
rect 350580 293724 350760 293812
rect 351014 293724 351194 293812
rect 351302 293724 351482 293812
rect 351590 293724 351770 293812
rect 351878 293724 352058 293812
rect 352166 293724 352346 293812
rect 352454 293724 352634 293812
rect 352742 293724 352922 293812
rect 353030 293724 353210 293812
rect 353464 293724 353644 293812
rect 353752 293724 353932 293812
rect 354040 293724 354220 293812
rect 354328 293724 354508 293812
rect 354616 293724 354796 293812
rect 354904 293724 355084 293812
rect 355192 293724 355372 293812
rect 355480 293724 355660 293812
rect 355914 293724 356094 293812
rect 356202 293724 356382 293812
rect 356490 293724 356670 293812
rect 356778 293724 356958 293812
rect 357066 293724 357246 293812
rect 357354 293724 357534 293812
rect 357642 293724 357822 293812
rect 357930 293724 358110 293812
rect 358364 293724 358544 293812
rect 358652 293724 358832 293812
rect 358940 293724 359120 293812
rect 359228 293724 359408 293812
rect 359516 293724 359696 293812
rect 359804 293724 359984 293812
rect 360092 293724 360272 293812
rect 360380 293724 360560 293812
rect 360814 293724 360994 293812
rect 361102 293724 361282 293812
rect 361390 293724 361570 293812
rect 361678 293724 361858 293812
rect 361966 293724 362146 293812
rect 362254 293724 362434 293812
rect 362542 293724 362722 293812
rect 362830 293724 363010 293812
rect 363264 293724 363444 293812
rect 363552 293724 363732 293812
rect 363840 293724 364020 293812
rect 364128 293724 364308 293812
rect 364416 293724 364596 293812
rect 364704 293724 364884 293812
rect 364992 293724 365172 293812
rect 365280 293724 365460 293812
rect 365714 293724 365894 293812
rect 366002 293724 366182 293812
rect 366290 293724 366470 293812
rect 366578 293724 366758 293812
rect 366866 293724 367046 293812
rect 367154 293724 367334 293812
rect 367442 293724 367622 293812
rect 367730 293724 367910 293812
rect 243214 293248 243394 293336
rect 243502 293248 243682 293336
rect 243790 293248 243970 293336
rect 244078 293248 244258 293336
rect 244366 293248 244546 293336
rect 244654 293248 244834 293336
rect 244942 293248 245122 293336
rect 245230 293248 245410 293336
rect 245664 293248 245844 293336
rect 245952 293248 246132 293336
rect 246240 293248 246420 293336
rect 246528 293248 246708 293336
rect 246816 293248 246996 293336
rect 247104 293248 247284 293336
rect 247392 293248 247572 293336
rect 247680 293248 247860 293336
rect 248114 293248 248294 293336
rect 248402 293248 248582 293336
rect 248690 293248 248870 293336
rect 248978 293248 249158 293336
rect 249266 293248 249446 293336
rect 249554 293248 249734 293336
rect 249842 293248 250022 293336
rect 250130 293248 250310 293336
rect 250564 293248 250744 293336
rect 250852 293248 251032 293336
rect 251140 293248 251320 293336
rect 251428 293248 251608 293336
rect 251716 293248 251896 293336
rect 252004 293248 252184 293336
rect 252292 293248 252472 293336
rect 252580 293248 252760 293336
rect 253014 293248 253194 293336
rect 253302 293248 253482 293336
rect 253590 293248 253770 293336
rect 253878 293248 254058 293336
rect 254166 293248 254346 293336
rect 254454 293248 254634 293336
rect 254742 293248 254922 293336
rect 255030 293248 255210 293336
rect 255464 293248 255644 293336
rect 255752 293248 255932 293336
rect 256040 293248 256220 293336
rect 256328 293248 256508 293336
rect 256616 293248 256796 293336
rect 256904 293248 257084 293336
rect 257192 293248 257372 293336
rect 257480 293248 257660 293336
rect 257914 293248 258094 293336
rect 258202 293248 258382 293336
rect 258490 293248 258670 293336
rect 258778 293248 258958 293336
rect 259066 293248 259246 293336
rect 259354 293248 259534 293336
rect 259642 293248 259822 293336
rect 259930 293248 260110 293336
rect 260364 293248 260544 293336
rect 260652 293248 260832 293336
rect 260940 293248 261120 293336
rect 261228 293248 261408 293336
rect 261516 293248 261696 293336
rect 261804 293248 261984 293336
rect 262092 293248 262272 293336
rect 262380 293248 262560 293336
rect 262814 293248 262994 293336
rect 263102 293248 263282 293336
rect 263390 293248 263570 293336
rect 263678 293248 263858 293336
rect 263966 293248 264146 293336
rect 264254 293248 264434 293336
rect 264542 293248 264722 293336
rect 264830 293248 265010 293336
rect 265264 293248 265444 293336
rect 265552 293248 265732 293336
rect 265840 293248 266020 293336
rect 266128 293248 266308 293336
rect 266416 293248 266596 293336
rect 266704 293248 266884 293336
rect 266992 293248 267172 293336
rect 267280 293248 267460 293336
rect 267714 293248 267894 293336
rect 268002 293248 268182 293336
rect 268290 293248 268470 293336
rect 268578 293248 268758 293336
rect 268866 293248 269046 293336
rect 269154 293248 269334 293336
rect 269442 293248 269622 293336
rect 269730 293248 269910 293336
rect 270164 293248 270344 293336
rect 270452 293248 270632 293336
rect 270740 293248 270920 293336
rect 271028 293248 271208 293336
rect 271316 293248 271496 293336
rect 271604 293248 271784 293336
rect 271892 293248 272072 293336
rect 272180 293248 272360 293336
rect 272614 293248 272794 293336
rect 272902 293248 273082 293336
rect 273190 293248 273370 293336
rect 273478 293248 273658 293336
rect 273766 293248 273946 293336
rect 274054 293248 274234 293336
rect 274342 293248 274522 293336
rect 274630 293248 274810 293336
rect 275064 293248 275244 293336
rect 275352 293248 275532 293336
rect 275640 293248 275820 293336
rect 275928 293248 276108 293336
rect 276216 293248 276396 293336
rect 276504 293248 276684 293336
rect 276792 293248 276972 293336
rect 277080 293248 277260 293336
rect 277514 293248 277694 293336
rect 277802 293248 277982 293336
rect 278090 293248 278270 293336
rect 278378 293248 278558 293336
rect 278666 293248 278846 293336
rect 278954 293248 279134 293336
rect 279242 293248 279422 293336
rect 279530 293248 279710 293336
rect 279964 293248 280144 293336
rect 280252 293248 280432 293336
rect 280540 293248 280720 293336
rect 280828 293248 281008 293336
rect 281116 293248 281296 293336
rect 281404 293248 281584 293336
rect 281692 293248 281872 293336
rect 281980 293248 282160 293336
rect 282414 293248 282594 293336
rect 282702 293248 282882 293336
rect 282990 293248 283170 293336
rect 283278 293248 283458 293336
rect 283566 293248 283746 293336
rect 283854 293248 284034 293336
rect 284142 293248 284322 293336
rect 284430 293248 284610 293336
rect 284864 293248 285044 293336
rect 285152 293248 285332 293336
rect 285440 293248 285620 293336
rect 285728 293248 285908 293336
rect 286016 293248 286196 293336
rect 286304 293248 286484 293336
rect 286592 293248 286772 293336
rect 286880 293248 287060 293336
rect 287314 293248 287494 293336
rect 287602 293248 287782 293336
rect 287890 293248 288070 293336
rect 288178 293248 288358 293336
rect 288466 293248 288646 293336
rect 288754 293248 288934 293336
rect 289042 293248 289222 293336
rect 289330 293248 289510 293336
rect 289764 293248 289944 293336
rect 290052 293248 290232 293336
rect 290340 293248 290520 293336
rect 290628 293248 290808 293336
rect 290916 293248 291096 293336
rect 291204 293248 291384 293336
rect 291492 293248 291672 293336
rect 291780 293248 291960 293336
rect 292214 293248 292394 293336
rect 292502 293248 292682 293336
rect 292790 293248 292970 293336
rect 293078 293248 293258 293336
rect 293366 293248 293546 293336
rect 293654 293248 293834 293336
rect 293942 293248 294122 293336
rect 294230 293248 294410 293336
rect 294664 293248 294844 293336
rect 294952 293248 295132 293336
rect 295240 293248 295420 293336
rect 295528 293248 295708 293336
rect 295816 293248 295996 293336
rect 296104 293248 296284 293336
rect 296392 293248 296572 293336
rect 296680 293248 296860 293336
rect 297114 293248 297294 293336
rect 297402 293248 297582 293336
rect 297690 293248 297870 293336
rect 297978 293248 298158 293336
rect 298266 293248 298446 293336
rect 298554 293248 298734 293336
rect 298842 293248 299022 293336
rect 299130 293248 299310 293336
rect 299564 293248 299744 293336
rect 299852 293248 300032 293336
rect 300140 293248 300320 293336
rect 300428 293248 300608 293336
rect 300716 293248 300896 293336
rect 301004 293248 301184 293336
rect 301292 293248 301472 293336
rect 301580 293248 301760 293336
rect 302014 293248 302194 293336
rect 302302 293248 302482 293336
rect 302590 293248 302770 293336
rect 302878 293248 303058 293336
rect 303166 293248 303346 293336
rect 303454 293248 303634 293336
rect 303742 293248 303922 293336
rect 304030 293248 304210 293336
rect 304464 293248 304644 293336
rect 304752 293248 304932 293336
rect 305040 293248 305220 293336
rect 305328 293248 305508 293336
rect 305616 293248 305796 293336
rect 305904 293248 306084 293336
rect 306192 293248 306372 293336
rect 306480 293248 306660 293336
rect 306914 293248 307094 293336
rect 307202 293248 307382 293336
rect 307490 293248 307670 293336
rect 307778 293248 307958 293336
rect 308066 293248 308246 293336
rect 308354 293248 308534 293336
rect 308642 293248 308822 293336
rect 308930 293248 309110 293336
rect 309364 293248 309544 293336
rect 309652 293248 309832 293336
rect 309940 293248 310120 293336
rect 310228 293248 310408 293336
rect 310516 293248 310696 293336
rect 310804 293248 310984 293336
rect 311092 293248 311272 293336
rect 311380 293248 311560 293336
rect 311814 293248 311994 293336
rect 312102 293248 312282 293336
rect 312390 293248 312570 293336
rect 312678 293248 312858 293336
rect 312966 293248 313146 293336
rect 313254 293248 313434 293336
rect 313542 293248 313722 293336
rect 313830 293248 314010 293336
rect 314264 293248 314444 293336
rect 314552 293248 314732 293336
rect 314840 293248 315020 293336
rect 315128 293248 315308 293336
rect 315416 293248 315596 293336
rect 315704 293248 315884 293336
rect 315992 293248 316172 293336
rect 316280 293248 316460 293336
rect 316714 293248 316894 293336
rect 317002 293248 317182 293336
rect 317290 293248 317470 293336
rect 317578 293248 317758 293336
rect 317866 293248 318046 293336
rect 318154 293248 318334 293336
rect 318442 293248 318622 293336
rect 318730 293248 318910 293336
rect 319164 293248 319344 293336
rect 319452 293248 319632 293336
rect 319740 293248 319920 293336
rect 320028 293248 320208 293336
rect 320316 293248 320496 293336
rect 320604 293248 320784 293336
rect 320892 293248 321072 293336
rect 321180 293248 321360 293336
rect 321614 293248 321794 293336
rect 321902 293248 322082 293336
rect 322190 293248 322370 293336
rect 322478 293248 322658 293336
rect 322766 293248 322946 293336
rect 323054 293248 323234 293336
rect 323342 293248 323522 293336
rect 323630 293248 323810 293336
rect 324064 293248 324244 293336
rect 324352 293248 324532 293336
rect 324640 293248 324820 293336
rect 324928 293248 325108 293336
rect 325216 293248 325396 293336
rect 325504 293248 325684 293336
rect 325792 293248 325972 293336
rect 326080 293248 326260 293336
rect 326514 293248 326694 293336
rect 326802 293248 326982 293336
rect 327090 293248 327270 293336
rect 327378 293248 327558 293336
rect 327666 293248 327846 293336
rect 327954 293248 328134 293336
rect 328242 293248 328422 293336
rect 328530 293248 328710 293336
rect 328964 293248 329144 293336
rect 329252 293248 329432 293336
rect 329540 293248 329720 293336
rect 329828 293248 330008 293336
rect 330116 293248 330296 293336
rect 330404 293248 330584 293336
rect 330692 293248 330872 293336
rect 330980 293248 331160 293336
rect 331414 293248 331594 293336
rect 331702 293248 331882 293336
rect 331990 293248 332170 293336
rect 332278 293248 332458 293336
rect 332566 293248 332746 293336
rect 332854 293248 333034 293336
rect 333142 293248 333322 293336
rect 333430 293248 333610 293336
rect 333864 293248 334044 293336
rect 334152 293248 334332 293336
rect 334440 293248 334620 293336
rect 334728 293248 334908 293336
rect 335016 293248 335196 293336
rect 335304 293248 335484 293336
rect 335592 293248 335772 293336
rect 335880 293248 336060 293336
rect 336314 293248 336494 293336
rect 336602 293248 336782 293336
rect 336890 293248 337070 293336
rect 337178 293248 337358 293336
rect 337466 293248 337646 293336
rect 337754 293248 337934 293336
rect 338042 293248 338222 293336
rect 338330 293248 338510 293336
rect 338764 293248 338944 293336
rect 339052 293248 339232 293336
rect 339340 293248 339520 293336
rect 339628 293248 339808 293336
rect 339916 293248 340096 293336
rect 340204 293248 340384 293336
rect 340492 293248 340672 293336
rect 340780 293248 340960 293336
rect 341214 293248 341394 293336
rect 341502 293248 341682 293336
rect 341790 293248 341970 293336
rect 342078 293248 342258 293336
rect 342366 293248 342546 293336
rect 342654 293248 342834 293336
rect 342942 293248 343122 293336
rect 343230 293248 343410 293336
rect 343664 293248 343844 293336
rect 343952 293248 344132 293336
rect 344240 293248 344420 293336
rect 344528 293248 344708 293336
rect 344816 293248 344996 293336
rect 345104 293248 345284 293336
rect 345392 293248 345572 293336
rect 345680 293248 345860 293336
rect 346114 293248 346294 293336
rect 346402 293248 346582 293336
rect 346690 293248 346870 293336
rect 346978 293248 347158 293336
rect 347266 293248 347446 293336
rect 347554 293248 347734 293336
rect 347842 293248 348022 293336
rect 348130 293248 348310 293336
rect 348564 293248 348744 293336
rect 348852 293248 349032 293336
rect 349140 293248 349320 293336
rect 349428 293248 349608 293336
rect 349716 293248 349896 293336
rect 350004 293248 350184 293336
rect 350292 293248 350472 293336
rect 350580 293248 350760 293336
rect 351014 293248 351194 293336
rect 351302 293248 351482 293336
rect 351590 293248 351770 293336
rect 351878 293248 352058 293336
rect 352166 293248 352346 293336
rect 352454 293248 352634 293336
rect 352742 293248 352922 293336
rect 353030 293248 353210 293336
rect 353464 293248 353644 293336
rect 353752 293248 353932 293336
rect 354040 293248 354220 293336
rect 354328 293248 354508 293336
rect 354616 293248 354796 293336
rect 354904 293248 355084 293336
rect 355192 293248 355372 293336
rect 355480 293248 355660 293336
rect 355914 293248 356094 293336
rect 356202 293248 356382 293336
rect 356490 293248 356670 293336
rect 356778 293248 356958 293336
rect 357066 293248 357246 293336
rect 357354 293248 357534 293336
rect 357642 293248 357822 293336
rect 357930 293248 358110 293336
rect 358364 293248 358544 293336
rect 358652 293248 358832 293336
rect 358940 293248 359120 293336
rect 359228 293248 359408 293336
rect 359516 293248 359696 293336
rect 359804 293248 359984 293336
rect 360092 293248 360272 293336
rect 360380 293248 360560 293336
rect 360814 293248 360994 293336
rect 361102 293248 361282 293336
rect 361390 293248 361570 293336
rect 361678 293248 361858 293336
rect 361966 293248 362146 293336
rect 362254 293248 362434 293336
rect 362542 293248 362722 293336
rect 362830 293248 363010 293336
rect 363264 293248 363444 293336
rect 363552 293248 363732 293336
rect 363840 293248 364020 293336
rect 364128 293248 364308 293336
rect 364416 293248 364596 293336
rect 364704 293248 364884 293336
rect 364992 293248 365172 293336
rect 365280 293248 365460 293336
rect 365714 293248 365894 293336
rect 366002 293248 366182 293336
rect 366290 293248 366470 293336
rect 366578 293248 366758 293336
rect 366866 293248 367046 293336
rect 367154 293248 367334 293336
rect 367442 293248 367622 293336
rect 367730 293248 367910 293336
rect 243214 293032 243394 293120
rect 243502 293032 243682 293120
rect 243790 293032 243970 293120
rect 244078 293032 244258 293120
rect 244366 293032 244546 293120
rect 244654 293032 244834 293120
rect 244942 293032 245122 293120
rect 245230 293032 245410 293120
rect 245664 293032 245844 293120
rect 245952 293032 246132 293120
rect 246240 293032 246420 293120
rect 246528 293032 246708 293120
rect 246816 293032 246996 293120
rect 247104 293032 247284 293120
rect 247392 293032 247572 293120
rect 247680 293032 247860 293120
rect 248114 293032 248294 293120
rect 248402 293032 248582 293120
rect 248690 293032 248870 293120
rect 248978 293032 249158 293120
rect 249266 293032 249446 293120
rect 249554 293032 249734 293120
rect 249842 293032 250022 293120
rect 250130 293032 250310 293120
rect 250564 293032 250744 293120
rect 250852 293032 251032 293120
rect 251140 293032 251320 293120
rect 251428 293032 251608 293120
rect 251716 293032 251896 293120
rect 252004 293032 252184 293120
rect 252292 293032 252472 293120
rect 252580 293032 252760 293120
rect 253014 293032 253194 293120
rect 253302 293032 253482 293120
rect 253590 293032 253770 293120
rect 253878 293032 254058 293120
rect 254166 293032 254346 293120
rect 254454 293032 254634 293120
rect 254742 293032 254922 293120
rect 255030 293032 255210 293120
rect 255464 293032 255644 293120
rect 255752 293032 255932 293120
rect 256040 293032 256220 293120
rect 256328 293032 256508 293120
rect 256616 293032 256796 293120
rect 256904 293032 257084 293120
rect 257192 293032 257372 293120
rect 257480 293032 257660 293120
rect 257914 293032 258094 293120
rect 258202 293032 258382 293120
rect 258490 293032 258670 293120
rect 258778 293032 258958 293120
rect 259066 293032 259246 293120
rect 259354 293032 259534 293120
rect 259642 293032 259822 293120
rect 259930 293032 260110 293120
rect 260364 293032 260544 293120
rect 260652 293032 260832 293120
rect 260940 293032 261120 293120
rect 261228 293032 261408 293120
rect 261516 293032 261696 293120
rect 261804 293032 261984 293120
rect 262092 293032 262272 293120
rect 262380 293032 262560 293120
rect 262814 293032 262994 293120
rect 263102 293032 263282 293120
rect 263390 293032 263570 293120
rect 263678 293032 263858 293120
rect 263966 293032 264146 293120
rect 264254 293032 264434 293120
rect 264542 293032 264722 293120
rect 264830 293032 265010 293120
rect 265264 293032 265444 293120
rect 265552 293032 265732 293120
rect 265840 293032 266020 293120
rect 266128 293032 266308 293120
rect 266416 293032 266596 293120
rect 266704 293032 266884 293120
rect 266992 293032 267172 293120
rect 267280 293032 267460 293120
rect 267714 293032 267894 293120
rect 268002 293032 268182 293120
rect 268290 293032 268470 293120
rect 268578 293032 268758 293120
rect 268866 293032 269046 293120
rect 269154 293032 269334 293120
rect 269442 293032 269622 293120
rect 269730 293032 269910 293120
rect 270164 293032 270344 293120
rect 270452 293032 270632 293120
rect 270740 293032 270920 293120
rect 271028 293032 271208 293120
rect 271316 293032 271496 293120
rect 271604 293032 271784 293120
rect 271892 293032 272072 293120
rect 272180 293032 272360 293120
rect 272614 293032 272794 293120
rect 272902 293032 273082 293120
rect 273190 293032 273370 293120
rect 273478 293032 273658 293120
rect 273766 293032 273946 293120
rect 274054 293032 274234 293120
rect 274342 293032 274522 293120
rect 274630 293032 274810 293120
rect 275064 293032 275244 293120
rect 275352 293032 275532 293120
rect 275640 293032 275820 293120
rect 275928 293032 276108 293120
rect 276216 293032 276396 293120
rect 276504 293032 276684 293120
rect 276792 293032 276972 293120
rect 277080 293032 277260 293120
rect 277514 293032 277694 293120
rect 277802 293032 277982 293120
rect 278090 293032 278270 293120
rect 278378 293032 278558 293120
rect 278666 293032 278846 293120
rect 278954 293032 279134 293120
rect 279242 293032 279422 293120
rect 279530 293032 279710 293120
rect 279964 293032 280144 293120
rect 280252 293032 280432 293120
rect 280540 293032 280720 293120
rect 280828 293032 281008 293120
rect 281116 293032 281296 293120
rect 281404 293032 281584 293120
rect 281692 293032 281872 293120
rect 281980 293032 282160 293120
rect 282414 293032 282594 293120
rect 282702 293032 282882 293120
rect 282990 293032 283170 293120
rect 283278 293032 283458 293120
rect 283566 293032 283746 293120
rect 283854 293032 284034 293120
rect 284142 293032 284322 293120
rect 284430 293032 284610 293120
rect 284864 293032 285044 293120
rect 285152 293032 285332 293120
rect 285440 293032 285620 293120
rect 285728 293032 285908 293120
rect 286016 293032 286196 293120
rect 286304 293032 286484 293120
rect 286592 293032 286772 293120
rect 286880 293032 287060 293120
rect 287314 293032 287494 293120
rect 287602 293032 287782 293120
rect 287890 293032 288070 293120
rect 288178 293032 288358 293120
rect 288466 293032 288646 293120
rect 288754 293032 288934 293120
rect 289042 293032 289222 293120
rect 289330 293032 289510 293120
rect 289764 293032 289944 293120
rect 290052 293032 290232 293120
rect 290340 293032 290520 293120
rect 290628 293032 290808 293120
rect 290916 293032 291096 293120
rect 291204 293032 291384 293120
rect 291492 293032 291672 293120
rect 291780 293032 291960 293120
rect 292214 293032 292394 293120
rect 292502 293032 292682 293120
rect 292790 293032 292970 293120
rect 293078 293032 293258 293120
rect 293366 293032 293546 293120
rect 293654 293032 293834 293120
rect 293942 293032 294122 293120
rect 294230 293032 294410 293120
rect 294664 293032 294844 293120
rect 294952 293032 295132 293120
rect 295240 293032 295420 293120
rect 295528 293032 295708 293120
rect 295816 293032 295996 293120
rect 296104 293032 296284 293120
rect 296392 293032 296572 293120
rect 296680 293032 296860 293120
rect 297114 293032 297294 293120
rect 297402 293032 297582 293120
rect 297690 293032 297870 293120
rect 297978 293032 298158 293120
rect 298266 293032 298446 293120
rect 298554 293032 298734 293120
rect 298842 293032 299022 293120
rect 299130 293032 299310 293120
rect 299564 293032 299744 293120
rect 299852 293032 300032 293120
rect 300140 293032 300320 293120
rect 300428 293032 300608 293120
rect 300716 293032 300896 293120
rect 301004 293032 301184 293120
rect 301292 293032 301472 293120
rect 301580 293032 301760 293120
rect 302014 293032 302194 293120
rect 302302 293032 302482 293120
rect 302590 293032 302770 293120
rect 302878 293032 303058 293120
rect 303166 293032 303346 293120
rect 303454 293032 303634 293120
rect 303742 293032 303922 293120
rect 304030 293032 304210 293120
rect 304464 293032 304644 293120
rect 304752 293032 304932 293120
rect 305040 293032 305220 293120
rect 305328 293032 305508 293120
rect 305616 293032 305796 293120
rect 305904 293032 306084 293120
rect 306192 293032 306372 293120
rect 306480 293032 306660 293120
rect 306914 293032 307094 293120
rect 307202 293032 307382 293120
rect 307490 293032 307670 293120
rect 307778 293032 307958 293120
rect 308066 293032 308246 293120
rect 308354 293032 308534 293120
rect 308642 293032 308822 293120
rect 308930 293032 309110 293120
rect 309364 293032 309544 293120
rect 309652 293032 309832 293120
rect 309940 293032 310120 293120
rect 310228 293032 310408 293120
rect 310516 293032 310696 293120
rect 310804 293032 310984 293120
rect 311092 293032 311272 293120
rect 311380 293032 311560 293120
rect 311814 293032 311994 293120
rect 312102 293032 312282 293120
rect 312390 293032 312570 293120
rect 312678 293032 312858 293120
rect 312966 293032 313146 293120
rect 313254 293032 313434 293120
rect 313542 293032 313722 293120
rect 313830 293032 314010 293120
rect 314264 293032 314444 293120
rect 314552 293032 314732 293120
rect 314840 293032 315020 293120
rect 315128 293032 315308 293120
rect 315416 293032 315596 293120
rect 315704 293032 315884 293120
rect 315992 293032 316172 293120
rect 316280 293032 316460 293120
rect 316714 293032 316894 293120
rect 317002 293032 317182 293120
rect 317290 293032 317470 293120
rect 317578 293032 317758 293120
rect 317866 293032 318046 293120
rect 318154 293032 318334 293120
rect 318442 293032 318622 293120
rect 318730 293032 318910 293120
rect 319164 293032 319344 293120
rect 319452 293032 319632 293120
rect 319740 293032 319920 293120
rect 320028 293032 320208 293120
rect 320316 293032 320496 293120
rect 320604 293032 320784 293120
rect 320892 293032 321072 293120
rect 321180 293032 321360 293120
rect 321614 293032 321794 293120
rect 321902 293032 322082 293120
rect 322190 293032 322370 293120
rect 322478 293032 322658 293120
rect 322766 293032 322946 293120
rect 323054 293032 323234 293120
rect 323342 293032 323522 293120
rect 323630 293032 323810 293120
rect 324064 293032 324244 293120
rect 324352 293032 324532 293120
rect 324640 293032 324820 293120
rect 324928 293032 325108 293120
rect 325216 293032 325396 293120
rect 325504 293032 325684 293120
rect 325792 293032 325972 293120
rect 326080 293032 326260 293120
rect 326514 293032 326694 293120
rect 326802 293032 326982 293120
rect 327090 293032 327270 293120
rect 327378 293032 327558 293120
rect 327666 293032 327846 293120
rect 327954 293032 328134 293120
rect 328242 293032 328422 293120
rect 328530 293032 328710 293120
rect 328964 293032 329144 293120
rect 329252 293032 329432 293120
rect 329540 293032 329720 293120
rect 329828 293032 330008 293120
rect 330116 293032 330296 293120
rect 330404 293032 330584 293120
rect 330692 293032 330872 293120
rect 330980 293032 331160 293120
rect 331414 293032 331594 293120
rect 331702 293032 331882 293120
rect 331990 293032 332170 293120
rect 332278 293032 332458 293120
rect 332566 293032 332746 293120
rect 332854 293032 333034 293120
rect 333142 293032 333322 293120
rect 333430 293032 333610 293120
rect 333864 293032 334044 293120
rect 334152 293032 334332 293120
rect 334440 293032 334620 293120
rect 334728 293032 334908 293120
rect 335016 293032 335196 293120
rect 335304 293032 335484 293120
rect 335592 293032 335772 293120
rect 335880 293032 336060 293120
rect 336314 293032 336494 293120
rect 336602 293032 336782 293120
rect 336890 293032 337070 293120
rect 337178 293032 337358 293120
rect 337466 293032 337646 293120
rect 337754 293032 337934 293120
rect 338042 293032 338222 293120
rect 338330 293032 338510 293120
rect 338764 293032 338944 293120
rect 339052 293032 339232 293120
rect 339340 293032 339520 293120
rect 339628 293032 339808 293120
rect 339916 293032 340096 293120
rect 340204 293032 340384 293120
rect 340492 293032 340672 293120
rect 340780 293032 340960 293120
rect 341214 293032 341394 293120
rect 341502 293032 341682 293120
rect 341790 293032 341970 293120
rect 342078 293032 342258 293120
rect 342366 293032 342546 293120
rect 342654 293032 342834 293120
rect 342942 293032 343122 293120
rect 343230 293032 343410 293120
rect 343664 293032 343844 293120
rect 343952 293032 344132 293120
rect 344240 293032 344420 293120
rect 344528 293032 344708 293120
rect 344816 293032 344996 293120
rect 345104 293032 345284 293120
rect 345392 293032 345572 293120
rect 345680 293032 345860 293120
rect 346114 293032 346294 293120
rect 346402 293032 346582 293120
rect 346690 293032 346870 293120
rect 346978 293032 347158 293120
rect 347266 293032 347446 293120
rect 347554 293032 347734 293120
rect 347842 293032 348022 293120
rect 348130 293032 348310 293120
rect 348564 293032 348744 293120
rect 348852 293032 349032 293120
rect 349140 293032 349320 293120
rect 349428 293032 349608 293120
rect 349716 293032 349896 293120
rect 350004 293032 350184 293120
rect 350292 293032 350472 293120
rect 350580 293032 350760 293120
rect 351014 293032 351194 293120
rect 351302 293032 351482 293120
rect 351590 293032 351770 293120
rect 351878 293032 352058 293120
rect 352166 293032 352346 293120
rect 352454 293032 352634 293120
rect 352742 293032 352922 293120
rect 353030 293032 353210 293120
rect 353464 293032 353644 293120
rect 353752 293032 353932 293120
rect 354040 293032 354220 293120
rect 354328 293032 354508 293120
rect 354616 293032 354796 293120
rect 354904 293032 355084 293120
rect 355192 293032 355372 293120
rect 355480 293032 355660 293120
rect 355914 293032 356094 293120
rect 356202 293032 356382 293120
rect 356490 293032 356670 293120
rect 356778 293032 356958 293120
rect 357066 293032 357246 293120
rect 357354 293032 357534 293120
rect 357642 293032 357822 293120
rect 357930 293032 358110 293120
rect 358364 293032 358544 293120
rect 358652 293032 358832 293120
rect 358940 293032 359120 293120
rect 359228 293032 359408 293120
rect 359516 293032 359696 293120
rect 359804 293032 359984 293120
rect 360092 293032 360272 293120
rect 360380 293032 360560 293120
rect 360814 293032 360994 293120
rect 361102 293032 361282 293120
rect 361390 293032 361570 293120
rect 361678 293032 361858 293120
rect 361966 293032 362146 293120
rect 362254 293032 362434 293120
rect 362542 293032 362722 293120
rect 362830 293032 363010 293120
rect 363264 293032 363444 293120
rect 363552 293032 363732 293120
rect 363840 293032 364020 293120
rect 364128 293032 364308 293120
rect 364416 293032 364596 293120
rect 364704 293032 364884 293120
rect 364992 293032 365172 293120
rect 365280 293032 365460 293120
rect 365714 293032 365894 293120
rect 366002 293032 366182 293120
rect 366290 293032 366470 293120
rect 366578 293032 366758 293120
rect 366866 293032 367046 293120
rect 367154 293032 367334 293120
rect 367442 293032 367622 293120
rect 367730 293032 367910 293120
rect 243214 292556 243394 292644
rect 243502 292556 243682 292644
rect 243790 292556 243970 292644
rect 244078 292556 244258 292644
rect 244366 292556 244546 292644
rect 244654 292556 244834 292644
rect 244942 292556 245122 292644
rect 245230 292556 245410 292644
rect 245664 292556 245844 292644
rect 245952 292556 246132 292644
rect 246240 292556 246420 292644
rect 246528 292556 246708 292644
rect 246816 292556 246996 292644
rect 247104 292556 247284 292644
rect 247392 292556 247572 292644
rect 247680 292556 247860 292644
rect 248114 292556 248294 292644
rect 248402 292556 248582 292644
rect 248690 292556 248870 292644
rect 248978 292556 249158 292644
rect 249266 292556 249446 292644
rect 249554 292556 249734 292644
rect 249842 292556 250022 292644
rect 250130 292556 250310 292644
rect 250564 292556 250744 292644
rect 250852 292556 251032 292644
rect 251140 292556 251320 292644
rect 251428 292556 251608 292644
rect 251716 292556 251896 292644
rect 252004 292556 252184 292644
rect 252292 292556 252472 292644
rect 252580 292556 252760 292644
rect 253014 292556 253194 292644
rect 253302 292556 253482 292644
rect 253590 292556 253770 292644
rect 253878 292556 254058 292644
rect 254166 292556 254346 292644
rect 254454 292556 254634 292644
rect 254742 292556 254922 292644
rect 255030 292556 255210 292644
rect 255464 292556 255644 292644
rect 255752 292556 255932 292644
rect 256040 292556 256220 292644
rect 256328 292556 256508 292644
rect 256616 292556 256796 292644
rect 256904 292556 257084 292644
rect 257192 292556 257372 292644
rect 257480 292556 257660 292644
rect 257914 292556 258094 292644
rect 258202 292556 258382 292644
rect 258490 292556 258670 292644
rect 258778 292556 258958 292644
rect 259066 292556 259246 292644
rect 259354 292556 259534 292644
rect 259642 292556 259822 292644
rect 259930 292556 260110 292644
rect 260364 292556 260544 292644
rect 260652 292556 260832 292644
rect 260940 292556 261120 292644
rect 261228 292556 261408 292644
rect 261516 292556 261696 292644
rect 261804 292556 261984 292644
rect 262092 292556 262272 292644
rect 262380 292556 262560 292644
rect 262814 292556 262994 292644
rect 263102 292556 263282 292644
rect 263390 292556 263570 292644
rect 263678 292556 263858 292644
rect 263966 292556 264146 292644
rect 264254 292556 264434 292644
rect 264542 292556 264722 292644
rect 264830 292556 265010 292644
rect 265264 292556 265444 292644
rect 265552 292556 265732 292644
rect 265840 292556 266020 292644
rect 266128 292556 266308 292644
rect 266416 292556 266596 292644
rect 266704 292556 266884 292644
rect 266992 292556 267172 292644
rect 267280 292556 267460 292644
rect 267714 292556 267894 292644
rect 268002 292556 268182 292644
rect 268290 292556 268470 292644
rect 268578 292556 268758 292644
rect 268866 292556 269046 292644
rect 269154 292556 269334 292644
rect 269442 292556 269622 292644
rect 269730 292556 269910 292644
rect 270164 292556 270344 292644
rect 270452 292556 270632 292644
rect 270740 292556 270920 292644
rect 271028 292556 271208 292644
rect 271316 292556 271496 292644
rect 271604 292556 271784 292644
rect 271892 292556 272072 292644
rect 272180 292556 272360 292644
rect 272614 292556 272794 292644
rect 272902 292556 273082 292644
rect 273190 292556 273370 292644
rect 273478 292556 273658 292644
rect 273766 292556 273946 292644
rect 274054 292556 274234 292644
rect 274342 292556 274522 292644
rect 274630 292556 274810 292644
rect 275064 292556 275244 292644
rect 275352 292556 275532 292644
rect 275640 292556 275820 292644
rect 275928 292556 276108 292644
rect 276216 292556 276396 292644
rect 276504 292556 276684 292644
rect 276792 292556 276972 292644
rect 277080 292556 277260 292644
rect 277514 292556 277694 292644
rect 277802 292556 277982 292644
rect 278090 292556 278270 292644
rect 278378 292556 278558 292644
rect 278666 292556 278846 292644
rect 278954 292556 279134 292644
rect 279242 292556 279422 292644
rect 279530 292556 279710 292644
rect 279964 292556 280144 292644
rect 280252 292556 280432 292644
rect 280540 292556 280720 292644
rect 280828 292556 281008 292644
rect 281116 292556 281296 292644
rect 281404 292556 281584 292644
rect 281692 292556 281872 292644
rect 281980 292556 282160 292644
rect 282414 292556 282594 292644
rect 282702 292556 282882 292644
rect 282990 292556 283170 292644
rect 283278 292556 283458 292644
rect 283566 292556 283746 292644
rect 283854 292556 284034 292644
rect 284142 292556 284322 292644
rect 284430 292556 284610 292644
rect 284864 292556 285044 292644
rect 285152 292556 285332 292644
rect 285440 292556 285620 292644
rect 285728 292556 285908 292644
rect 286016 292556 286196 292644
rect 286304 292556 286484 292644
rect 286592 292556 286772 292644
rect 286880 292556 287060 292644
rect 287314 292556 287494 292644
rect 287602 292556 287782 292644
rect 287890 292556 288070 292644
rect 288178 292556 288358 292644
rect 288466 292556 288646 292644
rect 288754 292556 288934 292644
rect 289042 292556 289222 292644
rect 289330 292556 289510 292644
rect 289764 292556 289944 292644
rect 290052 292556 290232 292644
rect 290340 292556 290520 292644
rect 290628 292556 290808 292644
rect 290916 292556 291096 292644
rect 291204 292556 291384 292644
rect 291492 292556 291672 292644
rect 291780 292556 291960 292644
rect 292214 292556 292394 292644
rect 292502 292556 292682 292644
rect 292790 292556 292970 292644
rect 293078 292556 293258 292644
rect 293366 292556 293546 292644
rect 293654 292556 293834 292644
rect 293942 292556 294122 292644
rect 294230 292556 294410 292644
rect 294664 292556 294844 292644
rect 294952 292556 295132 292644
rect 295240 292556 295420 292644
rect 295528 292556 295708 292644
rect 295816 292556 295996 292644
rect 296104 292556 296284 292644
rect 296392 292556 296572 292644
rect 296680 292556 296860 292644
rect 297114 292556 297294 292644
rect 297402 292556 297582 292644
rect 297690 292556 297870 292644
rect 297978 292556 298158 292644
rect 298266 292556 298446 292644
rect 298554 292556 298734 292644
rect 298842 292556 299022 292644
rect 299130 292556 299310 292644
rect 299564 292556 299744 292644
rect 299852 292556 300032 292644
rect 300140 292556 300320 292644
rect 300428 292556 300608 292644
rect 300716 292556 300896 292644
rect 301004 292556 301184 292644
rect 301292 292556 301472 292644
rect 301580 292556 301760 292644
rect 302014 292556 302194 292644
rect 302302 292556 302482 292644
rect 302590 292556 302770 292644
rect 302878 292556 303058 292644
rect 303166 292556 303346 292644
rect 303454 292556 303634 292644
rect 303742 292556 303922 292644
rect 304030 292556 304210 292644
rect 304464 292556 304644 292644
rect 304752 292556 304932 292644
rect 305040 292556 305220 292644
rect 305328 292556 305508 292644
rect 305616 292556 305796 292644
rect 305904 292556 306084 292644
rect 306192 292556 306372 292644
rect 306480 292556 306660 292644
rect 306914 292556 307094 292644
rect 307202 292556 307382 292644
rect 307490 292556 307670 292644
rect 307778 292556 307958 292644
rect 308066 292556 308246 292644
rect 308354 292556 308534 292644
rect 308642 292556 308822 292644
rect 308930 292556 309110 292644
rect 309364 292556 309544 292644
rect 309652 292556 309832 292644
rect 309940 292556 310120 292644
rect 310228 292556 310408 292644
rect 310516 292556 310696 292644
rect 310804 292556 310984 292644
rect 311092 292556 311272 292644
rect 311380 292556 311560 292644
rect 311814 292556 311994 292644
rect 312102 292556 312282 292644
rect 312390 292556 312570 292644
rect 312678 292556 312858 292644
rect 312966 292556 313146 292644
rect 313254 292556 313434 292644
rect 313542 292556 313722 292644
rect 313830 292556 314010 292644
rect 314264 292556 314444 292644
rect 314552 292556 314732 292644
rect 314840 292556 315020 292644
rect 315128 292556 315308 292644
rect 315416 292556 315596 292644
rect 315704 292556 315884 292644
rect 315992 292556 316172 292644
rect 316280 292556 316460 292644
rect 316714 292556 316894 292644
rect 317002 292556 317182 292644
rect 317290 292556 317470 292644
rect 317578 292556 317758 292644
rect 317866 292556 318046 292644
rect 318154 292556 318334 292644
rect 318442 292556 318622 292644
rect 318730 292556 318910 292644
rect 319164 292556 319344 292644
rect 319452 292556 319632 292644
rect 319740 292556 319920 292644
rect 320028 292556 320208 292644
rect 320316 292556 320496 292644
rect 320604 292556 320784 292644
rect 320892 292556 321072 292644
rect 321180 292556 321360 292644
rect 321614 292556 321794 292644
rect 321902 292556 322082 292644
rect 322190 292556 322370 292644
rect 322478 292556 322658 292644
rect 322766 292556 322946 292644
rect 323054 292556 323234 292644
rect 323342 292556 323522 292644
rect 323630 292556 323810 292644
rect 324064 292556 324244 292644
rect 324352 292556 324532 292644
rect 324640 292556 324820 292644
rect 324928 292556 325108 292644
rect 325216 292556 325396 292644
rect 325504 292556 325684 292644
rect 325792 292556 325972 292644
rect 326080 292556 326260 292644
rect 326514 292556 326694 292644
rect 326802 292556 326982 292644
rect 327090 292556 327270 292644
rect 327378 292556 327558 292644
rect 327666 292556 327846 292644
rect 327954 292556 328134 292644
rect 328242 292556 328422 292644
rect 328530 292556 328710 292644
rect 328964 292556 329144 292644
rect 329252 292556 329432 292644
rect 329540 292556 329720 292644
rect 329828 292556 330008 292644
rect 330116 292556 330296 292644
rect 330404 292556 330584 292644
rect 330692 292556 330872 292644
rect 330980 292556 331160 292644
rect 331414 292556 331594 292644
rect 331702 292556 331882 292644
rect 331990 292556 332170 292644
rect 332278 292556 332458 292644
rect 332566 292556 332746 292644
rect 332854 292556 333034 292644
rect 333142 292556 333322 292644
rect 333430 292556 333610 292644
rect 333864 292556 334044 292644
rect 334152 292556 334332 292644
rect 334440 292556 334620 292644
rect 334728 292556 334908 292644
rect 335016 292556 335196 292644
rect 335304 292556 335484 292644
rect 335592 292556 335772 292644
rect 335880 292556 336060 292644
rect 336314 292556 336494 292644
rect 336602 292556 336782 292644
rect 336890 292556 337070 292644
rect 337178 292556 337358 292644
rect 337466 292556 337646 292644
rect 337754 292556 337934 292644
rect 338042 292556 338222 292644
rect 338330 292556 338510 292644
rect 338764 292556 338944 292644
rect 339052 292556 339232 292644
rect 339340 292556 339520 292644
rect 339628 292556 339808 292644
rect 339916 292556 340096 292644
rect 340204 292556 340384 292644
rect 340492 292556 340672 292644
rect 340780 292556 340960 292644
rect 341214 292556 341394 292644
rect 341502 292556 341682 292644
rect 341790 292556 341970 292644
rect 342078 292556 342258 292644
rect 342366 292556 342546 292644
rect 342654 292556 342834 292644
rect 342942 292556 343122 292644
rect 343230 292556 343410 292644
rect 343664 292556 343844 292644
rect 343952 292556 344132 292644
rect 344240 292556 344420 292644
rect 344528 292556 344708 292644
rect 344816 292556 344996 292644
rect 345104 292556 345284 292644
rect 345392 292556 345572 292644
rect 345680 292556 345860 292644
rect 346114 292556 346294 292644
rect 346402 292556 346582 292644
rect 346690 292556 346870 292644
rect 346978 292556 347158 292644
rect 347266 292556 347446 292644
rect 347554 292556 347734 292644
rect 347842 292556 348022 292644
rect 348130 292556 348310 292644
rect 348564 292556 348744 292644
rect 348852 292556 349032 292644
rect 349140 292556 349320 292644
rect 349428 292556 349608 292644
rect 349716 292556 349896 292644
rect 350004 292556 350184 292644
rect 350292 292556 350472 292644
rect 350580 292556 350760 292644
rect 351014 292556 351194 292644
rect 351302 292556 351482 292644
rect 351590 292556 351770 292644
rect 351878 292556 352058 292644
rect 352166 292556 352346 292644
rect 352454 292556 352634 292644
rect 352742 292556 352922 292644
rect 353030 292556 353210 292644
rect 353464 292556 353644 292644
rect 353752 292556 353932 292644
rect 354040 292556 354220 292644
rect 354328 292556 354508 292644
rect 354616 292556 354796 292644
rect 354904 292556 355084 292644
rect 355192 292556 355372 292644
rect 355480 292556 355660 292644
rect 355914 292556 356094 292644
rect 356202 292556 356382 292644
rect 356490 292556 356670 292644
rect 356778 292556 356958 292644
rect 357066 292556 357246 292644
rect 357354 292556 357534 292644
rect 357642 292556 357822 292644
rect 357930 292556 358110 292644
rect 358364 292556 358544 292644
rect 358652 292556 358832 292644
rect 358940 292556 359120 292644
rect 359228 292556 359408 292644
rect 359516 292556 359696 292644
rect 359804 292556 359984 292644
rect 360092 292556 360272 292644
rect 360380 292556 360560 292644
rect 360814 292556 360994 292644
rect 361102 292556 361282 292644
rect 361390 292556 361570 292644
rect 361678 292556 361858 292644
rect 361966 292556 362146 292644
rect 362254 292556 362434 292644
rect 362542 292556 362722 292644
rect 362830 292556 363010 292644
rect 363264 292556 363444 292644
rect 363552 292556 363732 292644
rect 363840 292556 364020 292644
rect 364128 292556 364308 292644
rect 364416 292556 364596 292644
rect 364704 292556 364884 292644
rect 364992 292556 365172 292644
rect 365280 292556 365460 292644
rect 365714 292556 365894 292644
rect 366002 292556 366182 292644
rect 366290 292556 366470 292644
rect 366578 292556 366758 292644
rect 366866 292556 367046 292644
rect 367154 292556 367334 292644
rect 367442 292556 367622 292644
rect 367730 292556 367910 292644
rect 243214 292340 243394 292428
rect 243502 292340 243682 292428
rect 243790 292340 243970 292428
rect 244078 292340 244258 292428
rect 244366 292340 244546 292428
rect 244654 292340 244834 292428
rect 244942 292340 245122 292428
rect 245230 292340 245410 292428
rect 245664 292340 245844 292428
rect 245952 292340 246132 292428
rect 246240 292340 246420 292428
rect 246528 292340 246708 292428
rect 246816 292340 246996 292428
rect 247104 292340 247284 292428
rect 247392 292340 247572 292428
rect 247680 292340 247860 292428
rect 248114 292340 248294 292428
rect 248402 292340 248582 292428
rect 248690 292340 248870 292428
rect 248978 292340 249158 292428
rect 249266 292340 249446 292428
rect 249554 292340 249734 292428
rect 249842 292340 250022 292428
rect 250130 292340 250310 292428
rect 250564 292340 250744 292428
rect 250852 292340 251032 292428
rect 251140 292340 251320 292428
rect 251428 292340 251608 292428
rect 251716 292340 251896 292428
rect 252004 292340 252184 292428
rect 252292 292340 252472 292428
rect 252580 292340 252760 292428
rect 253014 292340 253194 292428
rect 253302 292340 253482 292428
rect 253590 292340 253770 292428
rect 253878 292340 254058 292428
rect 254166 292340 254346 292428
rect 254454 292340 254634 292428
rect 254742 292340 254922 292428
rect 255030 292340 255210 292428
rect 255464 292340 255644 292428
rect 255752 292340 255932 292428
rect 256040 292340 256220 292428
rect 256328 292340 256508 292428
rect 256616 292340 256796 292428
rect 256904 292340 257084 292428
rect 257192 292340 257372 292428
rect 257480 292340 257660 292428
rect 257914 292340 258094 292428
rect 258202 292340 258382 292428
rect 258490 292340 258670 292428
rect 258778 292340 258958 292428
rect 259066 292340 259246 292428
rect 259354 292340 259534 292428
rect 259642 292340 259822 292428
rect 259930 292340 260110 292428
rect 260364 292340 260544 292428
rect 260652 292340 260832 292428
rect 260940 292340 261120 292428
rect 261228 292340 261408 292428
rect 261516 292340 261696 292428
rect 261804 292340 261984 292428
rect 262092 292340 262272 292428
rect 262380 292340 262560 292428
rect 262814 292340 262994 292428
rect 263102 292340 263282 292428
rect 263390 292340 263570 292428
rect 263678 292340 263858 292428
rect 263966 292340 264146 292428
rect 264254 292340 264434 292428
rect 264542 292340 264722 292428
rect 264830 292340 265010 292428
rect 265264 292340 265444 292428
rect 265552 292340 265732 292428
rect 265840 292340 266020 292428
rect 266128 292340 266308 292428
rect 266416 292340 266596 292428
rect 266704 292340 266884 292428
rect 266992 292340 267172 292428
rect 267280 292340 267460 292428
rect 267714 292340 267894 292428
rect 268002 292340 268182 292428
rect 268290 292340 268470 292428
rect 268578 292340 268758 292428
rect 268866 292340 269046 292428
rect 269154 292340 269334 292428
rect 269442 292340 269622 292428
rect 269730 292340 269910 292428
rect 270164 292340 270344 292428
rect 270452 292340 270632 292428
rect 270740 292340 270920 292428
rect 271028 292340 271208 292428
rect 271316 292340 271496 292428
rect 271604 292340 271784 292428
rect 271892 292340 272072 292428
rect 272180 292340 272360 292428
rect 272614 292340 272794 292428
rect 272902 292340 273082 292428
rect 273190 292340 273370 292428
rect 273478 292340 273658 292428
rect 273766 292340 273946 292428
rect 274054 292340 274234 292428
rect 274342 292340 274522 292428
rect 274630 292340 274810 292428
rect 275064 292340 275244 292428
rect 275352 292340 275532 292428
rect 275640 292340 275820 292428
rect 275928 292340 276108 292428
rect 276216 292340 276396 292428
rect 276504 292340 276684 292428
rect 276792 292340 276972 292428
rect 277080 292340 277260 292428
rect 277514 292340 277694 292428
rect 277802 292340 277982 292428
rect 278090 292340 278270 292428
rect 278378 292340 278558 292428
rect 278666 292340 278846 292428
rect 278954 292340 279134 292428
rect 279242 292340 279422 292428
rect 279530 292340 279710 292428
rect 279964 292340 280144 292428
rect 280252 292340 280432 292428
rect 280540 292340 280720 292428
rect 280828 292340 281008 292428
rect 281116 292340 281296 292428
rect 281404 292340 281584 292428
rect 281692 292340 281872 292428
rect 281980 292340 282160 292428
rect 282414 292340 282594 292428
rect 282702 292340 282882 292428
rect 282990 292340 283170 292428
rect 283278 292340 283458 292428
rect 283566 292340 283746 292428
rect 283854 292340 284034 292428
rect 284142 292340 284322 292428
rect 284430 292340 284610 292428
rect 284864 292340 285044 292428
rect 285152 292340 285332 292428
rect 285440 292340 285620 292428
rect 285728 292340 285908 292428
rect 286016 292340 286196 292428
rect 286304 292340 286484 292428
rect 286592 292340 286772 292428
rect 286880 292340 287060 292428
rect 287314 292340 287494 292428
rect 287602 292340 287782 292428
rect 287890 292340 288070 292428
rect 288178 292340 288358 292428
rect 288466 292340 288646 292428
rect 288754 292340 288934 292428
rect 289042 292340 289222 292428
rect 289330 292340 289510 292428
rect 289764 292340 289944 292428
rect 290052 292340 290232 292428
rect 290340 292340 290520 292428
rect 290628 292340 290808 292428
rect 290916 292340 291096 292428
rect 291204 292340 291384 292428
rect 291492 292340 291672 292428
rect 291780 292340 291960 292428
rect 292214 292340 292394 292428
rect 292502 292340 292682 292428
rect 292790 292340 292970 292428
rect 293078 292340 293258 292428
rect 293366 292340 293546 292428
rect 293654 292340 293834 292428
rect 293942 292340 294122 292428
rect 294230 292340 294410 292428
rect 294664 292340 294844 292428
rect 294952 292340 295132 292428
rect 295240 292340 295420 292428
rect 295528 292340 295708 292428
rect 295816 292340 295996 292428
rect 296104 292340 296284 292428
rect 296392 292340 296572 292428
rect 296680 292340 296860 292428
rect 297114 292340 297294 292428
rect 297402 292340 297582 292428
rect 297690 292340 297870 292428
rect 297978 292340 298158 292428
rect 298266 292340 298446 292428
rect 298554 292340 298734 292428
rect 298842 292340 299022 292428
rect 299130 292340 299310 292428
rect 299564 292340 299744 292428
rect 299852 292340 300032 292428
rect 300140 292340 300320 292428
rect 300428 292340 300608 292428
rect 300716 292340 300896 292428
rect 301004 292340 301184 292428
rect 301292 292340 301472 292428
rect 301580 292340 301760 292428
rect 302014 292340 302194 292428
rect 302302 292340 302482 292428
rect 302590 292340 302770 292428
rect 302878 292340 303058 292428
rect 303166 292340 303346 292428
rect 303454 292340 303634 292428
rect 303742 292340 303922 292428
rect 304030 292340 304210 292428
rect 304464 292340 304644 292428
rect 304752 292340 304932 292428
rect 305040 292340 305220 292428
rect 305328 292340 305508 292428
rect 305616 292340 305796 292428
rect 305904 292340 306084 292428
rect 306192 292340 306372 292428
rect 306480 292340 306660 292428
rect 306914 292340 307094 292428
rect 307202 292340 307382 292428
rect 307490 292340 307670 292428
rect 307778 292340 307958 292428
rect 308066 292340 308246 292428
rect 308354 292340 308534 292428
rect 308642 292340 308822 292428
rect 308930 292340 309110 292428
rect 309364 292340 309544 292428
rect 309652 292340 309832 292428
rect 309940 292340 310120 292428
rect 310228 292340 310408 292428
rect 310516 292340 310696 292428
rect 310804 292340 310984 292428
rect 311092 292340 311272 292428
rect 311380 292340 311560 292428
rect 311814 292340 311994 292428
rect 312102 292340 312282 292428
rect 312390 292340 312570 292428
rect 312678 292340 312858 292428
rect 312966 292340 313146 292428
rect 313254 292340 313434 292428
rect 313542 292340 313722 292428
rect 313830 292340 314010 292428
rect 314264 292340 314444 292428
rect 314552 292340 314732 292428
rect 314840 292340 315020 292428
rect 315128 292340 315308 292428
rect 315416 292340 315596 292428
rect 315704 292340 315884 292428
rect 315992 292340 316172 292428
rect 316280 292340 316460 292428
rect 316714 292340 316894 292428
rect 317002 292340 317182 292428
rect 317290 292340 317470 292428
rect 317578 292340 317758 292428
rect 317866 292340 318046 292428
rect 318154 292340 318334 292428
rect 318442 292340 318622 292428
rect 318730 292340 318910 292428
rect 319164 292340 319344 292428
rect 319452 292340 319632 292428
rect 319740 292340 319920 292428
rect 320028 292340 320208 292428
rect 320316 292340 320496 292428
rect 320604 292340 320784 292428
rect 320892 292340 321072 292428
rect 321180 292340 321360 292428
rect 321614 292340 321794 292428
rect 321902 292340 322082 292428
rect 322190 292340 322370 292428
rect 322478 292340 322658 292428
rect 322766 292340 322946 292428
rect 323054 292340 323234 292428
rect 323342 292340 323522 292428
rect 323630 292340 323810 292428
rect 324064 292340 324244 292428
rect 324352 292340 324532 292428
rect 324640 292340 324820 292428
rect 324928 292340 325108 292428
rect 325216 292340 325396 292428
rect 325504 292340 325684 292428
rect 325792 292340 325972 292428
rect 326080 292340 326260 292428
rect 326514 292340 326694 292428
rect 326802 292340 326982 292428
rect 327090 292340 327270 292428
rect 327378 292340 327558 292428
rect 327666 292340 327846 292428
rect 327954 292340 328134 292428
rect 328242 292340 328422 292428
rect 328530 292340 328710 292428
rect 328964 292340 329144 292428
rect 329252 292340 329432 292428
rect 329540 292340 329720 292428
rect 329828 292340 330008 292428
rect 330116 292340 330296 292428
rect 330404 292340 330584 292428
rect 330692 292340 330872 292428
rect 330980 292340 331160 292428
rect 331414 292340 331594 292428
rect 331702 292340 331882 292428
rect 331990 292340 332170 292428
rect 332278 292340 332458 292428
rect 332566 292340 332746 292428
rect 332854 292340 333034 292428
rect 333142 292340 333322 292428
rect 333430 292340 333610 292428
rect 333864 292340 334044 292428
rect 334152 292340 334332 292428
rect 334440 292340 334620 292428
rect 334728 292340 334908 292428
rect 335016 292340 335196 292428
rect 335304 292340 335484 292428
rect 335592 292340 335772 292428
rect 335880 292340 336060 292428
rect 336314 292340 336494 292428
rect 336602 292340 336782 292428
rect 336890 292340 337070 292428
rect 337178 292340 337358 292428
rect 337466 292340 337646 292428
rect 337754 292340 337934 292428
rect 338042 292340 338222 292428
rect 338330 292340 338510 292428
rect 338764 292340 338944 292428
rect 339052 292340 339232 292428
rect 339340 292340 339520 292428
rect 339628 292340 339808 292428
rect 339916 292340 340096 292428
rect 340204 292340 340384 292428
rect 340492 292340 340672 292428
rect 340780 292340 340960 292428
rect 341214 292340 341394 292428
rect 341502 292340 341682 292428
rect 341790 292340 341970 292428
rect 342078 292340 342258 292428
rect 342366 292340 342546 292428
rect 342654 292340 342834 292428
rect 342942 292340 343122 292428
rect 343230 292340 343410 292428
rect 343664 292340 343844 292428
rect 343952 292340 344132 292428
rect 344240 292340 344420 292428
rect 344528 292340 344708 292428
rect 344816 292340 344996 292428
rect 345104 292340 345284 292428
rect 345392 292340 345572 292428
rect 345680 292340 345860 292428
rect 346114 292340 346294 292428
rect 346402 292340 346582 292428
rect 346690 292340 346870 292428
rect 346978 292340 347158 292428
rect 347266 292340 347446 292428
rect 347554 292340 347734 292428
rect 347842 292340 348022 292428
rect 348130 292340 348310 292428
rect 348564 292340 348744 292428
rect 348852 292340 349032 292428
rect 349140 292340 349320 292428
rect 349428 292340 349608 292428
rect 349716 292340 349896 292428
rect 350004 292340 350184 292428
rect 350292 292340 350472 292428
rect 350580 292340 350760 292428
rect 351014 292340 351194 292428
rect 351302 292340 351482 292428
rect 351590 292340 351770 292428
rect 351878 292340 352058 292428
rect 352166 292340 352346 292428
rect 352454 292340 352634 292428
rect 352742 292340 352922 292428
rect 353030 292340 353210 292428
rect 353464 292340 353644 292428
rect 353752 292340 353932 292428
rect 354040 292340 354220 292428
rect 354328 292340 354508 292428
rect 354616 292340 354796 292428
rect 354904 292340 355084 292428
rect 355192 292340 355372 292428
rect 355480 292340 355660 292428
rect 355914 292340 356094 292428
rect 356202 292340 356382 292428
rect 356490 292340 356670 292428
rect 356778 292340 356958 292428
rect 357066 292340 357246 292428
rect 357354 292340 357534 292428
rect 357642 292340 357822 292428
rect 357930 292340 358110 292428
rect 358364 292340 358544 292428
rect 358652 292340 358832 292428
rect 358940 292340 359120 292428
rect 359228 292340 359408 292428
rect 359516 292340 359696 292428
rect 359804 292340 359984 292428
rect 360092 292340 360272 292428
rect 360380 292340 360560 292428
rect 360814 292340 360994 292428
rect 361102 292340 361282 292428
rect 361390 292340 361570 292428
rect 361678 292340 361858 292428
rect 361966 292340 362146 292428
rect 362254 292340 362434 292428
rect 362542 292340 362722 292428
rect 362830 292340 363010 292428
rect 363264 292340 363444 292428
rect 363552 292340 363732 292428
rect 363840 292340 364020 292428
rect 364128 292340 364308 292428
rect 364416 292340 364596 292428
rect 364704 292340 364884 292428
rect 364992 292340 365172 292428
rect 365280 292340 365460 292428
rect 365714 292340 365894 292428
rect 366002 292340 366182 292428
rect 366290 292340 366470 292428
rect 366578 292340 366758 292428
rect 366866 292340 367046 292428
rect 367154 292340 367334 292428
rect 367442 292340 367622 292428
rect 367730 292340 367910 292428
rect 243214 291864 243394 291952
rect 243502 291864 243682 291952
rect 243790 291864 243970 291952
rect 244078 291864 244258 291952
rect 244366 291864 244546 291952
rect 244654 291864 244834 291952
rect 244942 291864 245122 291952
rect 245230 291864 245410 291952
rect 245664 291864 245844 291952
rect 245952 291864 246132 291952
rect 246240 291864 246420 291952
rect 246528 291864 246708 291952
rect 246816 291864 246996 291952
rect 247104 291864 247284 291952
rect 247392 291864 247572 291952
rect 247680 291864 247860 291952
rect 248114 291864 248294 291952
rect 248402 291864 248582 291952
rect 248690 291864 248870 291952
rect 248978 291864 249158 291952
rect 249266 291864 249446 291952
rect 249554 291864 249734 291952
rect 249842 291864 250022 291952
rect 250130 291864 250310 291952
rect 250564 291864 250744 291952
rect 250852 291864 251032 291952
rect 251140 291864 251320 291952
rect 251428 291864 251608 291952
rect 251716 291864 251896 291952
rect 252004 291864 252184 291952
rect 252292 291864 252472 291952
rect 252580 291864 252760 291952
rect 253014 291864 253194 291952
rect 253302 291864 253482 291952
rect 253590 291864 253770 291952
rect 253878 291864 254058 291952
rect 254166 291864 254346 291952
rect 254454 291864 254634 291952
rect 254742 291864 254922 291952
rect 255030 291864 255210 291952
rect 255464 291864 255644 291952
rect 255752 291864 255932 291952
rect 256040 291864 256220 291952
rect 256328 291864 256508 291952
rect 256616 291864 256796 291952
rect 256904 291864 257084 291952
rect 257192 291864 257372 291952
rect 257480 291864 257660 291952
rect 257914 291864 258094 291952
rect 258202 291864 258382 291952
rect 258490 291864 258670 291952
rect 258778 291864 258958 291952
rect 259066 291864 259246 291952
rect 259354 291864 259534 291952
rect 259642 291864 259822 291952
rect 259930 291864 260110 291952
rect 260364 291864 260544 291952
rect 260652 291864 260832 291952
rect 260940 291864 261120 291952
rect 261228 291864 261408 291952
rect 261516 291864 261696 291952
rect 261804 291864 261984 291952
rect 262092 291864 262272 291952
rect 262380 291864 262560 291952
rect 262814 291864 262994 291952
rect 263102 291864 263282 291952
rect 263390 291864 263570 291952
rect 263678 291864 263858 291952
rect 263966 291864 264146 291952
rect 264254 291864 264434 291952
rect 264542 291864 264722 291952
rect 264830 291864 265010 291952
rect 265264 291864 265444 291952
rect 265552 291864 265732 291952
rect 265840 291864 266020 291952
rect 266128 291864 266308 291952
rect 266416 291864 266596 291952
rect 266704 291864 266884 291952
rect 266992 291864 267172 291952
rect 267280 291864 267460 291952
rect 267714 291864 267894 291952
rect 268002 291864 268182 291952
rect 268290 291864 268470 291952
rect 268578 291864 268758 291952
rect 268866 291864 269046 291952
rect 269154 291864 269334 291952
rect 269442 291864 269622 291952
rect 269730 291864 269910 291952
rect 270164 291864 270344 291952
rect 270452 291864 270632 291952
rect 270740 291864 270920 291952
rect 271028 291864 271208 291952
rect 271316 291864 271496 291952
rect 271604 291864 271784 291952
rect 271892 291864 272072 291952
rect 272180 291864 272360 291952
rect 272614 291864 272794 291952
rect 272902 291864 273082 291952
rect 273190 291864 273370 291952
rect 273478 291864 273658 291952
rect 273766 291864 273946 291952
rect 274054 291864 274234 291952
rect 274342 291864 274522 291952
rect 274630 291864 274810 291952
rect 275064 291864 275244 291952
rect 275352 291864 275532 291952
rect 275640 291864 275820 291952
rect 275928 291864 276108 291952
rect 276216 291864 276396 291952
rect 276504 291864 276684 291952
rect 276792 291864 276972 291952
rect 277080 291864 277260 291952
rect 277514 291864 277694 291952
rect 277802 291864 277982 291952
rect 278090 291864 278270 291952
rect 278378 291864 278558 291952
rect 278666 291864 278846 291952
rect 278954 291864 279134 291952
rect 279242 291864 279422 291952
rect 279530 291864 279710 291952
rect 279964 291864 280144 291952
rect 280252 291864 280432 291952
rect 280540 291864 280720 291952
rect 280828 291864 281008 291952
rect 281116 291864 281296 291952
rect 281404 291864 281584 291952
rect 281692 291864 281872 291952
rect 281980 291864 282160 291952
rect 282414 291864 282594 291952
rect 282702 291864 282882 291952
rect 282990 291864 283170 291952
rect 283278 291864 283458 291952
rect 283566 291864 283746 291952
rect 283854 291864 284034 291952
rect 284142 291864 284322 291952
rect 284430 291864 284610 291952
rect 284864 291864 285044 291952
rect 285152 291864 285332 291952
rect 285440 291864 285620 291952
rect 285728 291864 285908 291952
rect 286016 291864 286196 291952
rect 286304 291864 286484 291952
rect 286592 291864 286772 291952
rect 286880 291864 287060 291952
rect 287314 291864 287494 291952
rect 287602 291864 287782 291952
rect 287890 291864 288070 291952
rect 288178 291864 288358 291952
rect 288466 291864 288646 291952
rect 288754 291864 288934 291952
rect 289042 291864 289222 291952
rect 289330 291864 289510 291952
rect 289764 291864 289944 291952
rect 290052 291864 290232 291952
rect 290340 291864 290520 291952
rect 290628 291864 290808 291952
rect 290916 291864 291096 291952
rect 291204 291864 291384 291952
rect 291492 291864 291672 291952
rect 291780 291864 291960 291952
rect 292214 291864 292394 291952
rect 292502 291864 292682 291952
rect 292790 291864 292970 291952
rect 293078 291864 293258 291952
rect 293366 291864 293546 291952
rect 293654 291864 293834 291952
rect 293942 291864 294122 291952
rect 294230 291864 294410 291952
rect 294664 291864 294844 291952
rect 294952 291864 295132 291952
rect 295240 291864 295420 291952
rect 295528 291864 295708 291952
rect 295816 291864 295996 291952
rect 296104 291864 296284 291952
rect 296392 291864 296572 291952
rect 296680 291864 296860 291952
rect 297114 291864 297294 291952
rect 297402 291864 297582 291952
rect 297690 291864 297870 291952
rect 297978 291864 298158 291952
rect 298266 291864 298446 291952
rect 298554 291864 298734 291952
rect 298842 291864 299022 291952
rect 299130 291864 299310 291952
rect 299564 291864 299744 291952
rect 299852 291864 300032 291952
rect 300140 291864 300320 291952
rect 300428 291864 300608 291952
rect 300716 291864 300896 291952
rect 301004 291864 301184 291952
rect 301292 291864 301472 291952
rect 301580 291864 301760 291952
rect 302014 291864 302194 291952
rect 302302 291864 302482 291952
rect 302590 291864 302770 291952
rect 302878 291864 303058 291952
rect 303166 291864 303346 291952
rect 303454 291864 303634 291952
rect 303742 291864 303922 291952
rect 304030 291864 304210 291952
rect 304464 291864 304644 291952
rect 304752 291864 304932 291952
rect 305040 291864 305220 291952
rect 305328 291864 305508 291952
rect 305616 291864 305796 291952
rect 305904 291864 306084 291952
rect 306192 291864 306372 291952
rect 306480 291864 306660 291952
rect 306914 291864 307094 291952
rect 307202 291864 307382 291952
rect 307490 291864 307670 291952
rect 307778 291864 307958 291952
rect 308066 291864 308246 291952
rect 308354 291864 308534 291952
rect 308642 291864 308822 291952
rect 308930 291864 309110 291952
rect 309364 291864 309544 291952
rect 309652 291864 309832 291952
rect 309940 291864 310120 291952
rect 310228 291864 310408 291952
rect 310516 291864 310696 291952
rect 310804 291864 310984 291952
rect 311092 291864 311272 291952
rect 311380 291864 311560 291952
rect 311814 291864 311994 291952
rect 312102 291864 312282 291952
rect 312390 291864 312570 291952
rect 312678 291864 312858 291952
rect 312966 291864 313146 291952
rect 313254 291864 313434 291952
rect 313542 291864 313722 291952
rect 313830 291864 314010 291952
rect 314264 291864 314444 291952
rect 314552 291864 314732 291952
rect 314840 291864 315020 291952
rect 315128 291864 315308 291952
rect 315416 291864 315596 291952
rect 315704 291864 315884 291952
rect 315992 291864 316172 291952
rect 316280 291864 316460 291952
rect 316714 291864 316894 291952
rect 317002 291864 317182 291952
rect 317290 291864 317470 291952
rect 317578 291864 317758 291952
rect 317866 291864 318046 291952
rect 318154 291864 318334 291952
rect 318442 291864 318622 291952
rect 318730 291864 318910 291952
rect 319164 291864 319344 291952
rect 319452 291864 319632 291952
rect 319740 291864 319920 291952
rect 320028 291864 320208 291952
rect 320316 291864 320496 291952
rect 320604 291864 320784 291952
rect 320892 291864 321072 291952
rect 321180 291864 321360 291952
rect 321614 291864 321794 291952
rect 321902 291864 322082 291952
rect 322190 291864 322370 291952
rect 322478 291864 322658 291952
rect 322766 291864 322946 291952
rect 323054 291864 323234 291952
rect 323342 291864 323522 291952
rect 323630 291864 323810 291952
rect 324064 291864 324244 291952
rect 324352 291864 324532 291952
rect 324640 291864 324820 291952
rect 324928 291864 325108 291952
rect 325216 291864 325396 291952
rect 325504 291864 325684 291952
rect 325792 291864 325972 291952
rect 326080 291864 326260 291952
rect 326514 291864 326694 291952
rect 326802 291864 326982 291952
rect 327090 291864 327270 291952
rect 327378 291864 327558 291952
rect 327666 291864 327846 291952
rect 327954 291864 328134 291952
rect 328242 291864 328422 291952
rect 328530 291864 328710 291952
rect 328964 291864 329144 291952
rect 329252 291864 329432 291952
rect 329540 291864 329720 291952
rect 329828 291864 330008 291952
rect 330116 291864 330296 291952
rect 330404 291864 330584 291952
rect 330692 291864 330872 291952
rect 330980 291864 331160 291952
rect 331414 291864 331594 291952
rect 331702 291864 331882 291952
rect 331990 291864 332170 291952
rect 332278 291864 332458 291952
rect 332566 291864 332746 291952
rect 332854 291864 333034 291952
rect 333142 291864 333322 291952
rect 333430 291864 333610 291952
rect 333864 291864 334044 291952
rect 334152 291864 334332 291952
rect 334440 291864 334620 291952
rect 334728 291864 334908 291952
rect 335016 291864 335196 291952
rect 335304 291864 335484 291952
rect 335592 291864 335772 291952
rect 335880 291864 336060 291952
rect 336314 291864 336494 291952
rect 336602 291864 336782 291952
rect 336890 291864 337070 291952
rect 337178 291864 337358 291952
rect 337466 291864 337646 291952
rect 337754 291864 337934 291952
rect 338042 291864 338222 291952
rect 338330 291864 338510 291952
rect 338764 291864 338944 291952
rect 339052 291864 339232 291952
rect 339340 291864 339520 291952
rect 339628 291864 339808 291952
rect 339916 291864 340096 291952
rect 340204 291864 340384 291952
rect 340492 291864 340672 291952
rect 340780 291864 340960 291952
rect 341214 291864 341394 291952
rect 341502 291864 341682 291952
rect 341790 291864 341970 291952
rect 342078 291864 342258 291952
rect 342366 291864 342546 291952
rect 342654 291864 342834 291952
rect 342942 291864 343122 291952
rect 343230 291864 343410 291952
rect 343664 291864 343844 291952
rect 343952 291864 344132 291952
rect 344240 291864 344420 291952
rect 344528 291864 344708 291952
rect 344816 291864 344996 291952
rect 345104 291864 345284 291952
rect 345392 291864 345572 291952
rect 345680 291864 345860 291952
rect 346114 291864 346294 291952
rect 346402 291864 346582 291952
rect 346690 291864 346870 291952
rect 346978 291864 347158 291952
rect 347266 291864 347446 291952
rect 347554 291864 347734 291952
rect 347842 291864 348022 291952
rect 348130 291864 348310 291952
rect 348564 291864 348744 291952
rect 348852 291864 349032 291952
rect 349140 291864 349320 291952
rect 349428 291864 349608 291952
rect 349716 291864 349896 291952
rect 350004 291864 350184 291952
rect 350292 291864 350472 291952
rect 350580 291864 350760 291952
rect 351014 291864 351194 291952
rect 351302 291864 351482 291952
rect 351590 291864 351770 291952
rect 351878 291864 352058 291952
rect 352166 291864 352346 291952
rect 352454 291864 352634 291952
rect 352742 291864 352922 291952
rect 353030 291864 353210 291952
rect 353464 291864 353644 291952
rect 353752 291864 353932 291952
rect 354040 291864 354220 291952
rect 354328 291864 354508 291952
rect 354616 291864 354796 291952
rect 354904 291864 355084 291952
rect 355192 291864 355372 291952
rect 355480 291864 355660 291952
rect 355914 291864 356094 291952
rect 356202 291864 356382 291952
rect 356490 291864 356670 291952
rect 356778 291864 356958 291952
rect 357066 291864 357246 291952
rect 357354 291864 357534 291952
rect 357642 291864 357822 291952
rect 357930 291864 358110 291952
rect 358364 291864 358544 291952
rect 358652 291864 358832 291952
rect 358940 291864 359120 291952
rect 359228 291864 359408 291952
rect 359516 291864 359696 291952
rect 359804 291864 359984 291952
rect 360092 291864 360272 291952
rect 360380 291864 360560 291952
rect 360814 291864 360994 291952
rect 361102 291864 361282 291952
rect 361390 291864 361570 291952
rect 361678 291864 361858 291952
rect 361966 291864 362146 291952
rect 362254 291864 362434 291952
rect 362542 291864 362722 291952
rect 362830 291864 363010 291952
rect 363264 291864 363444 291952
rect 363552 291864 363732 291952
rect 363840 291864 364020 291952
rect 364128 291864 364308 291952
rect 364416 291864 364596 291952
rect 364704 291864 364884 291952
rect 364992 291864 365172 291952
rect 365280 291864 365460 291952
rect 365714 291864 365894 291952
rect 366002 291864 366182 291952
rect 366290 291864 366470 291952
rect 366578 291864 366758 291952
rect 366866 291864 367046 291952
rect 367154 291864 367334 291952
rect 367442 291864 367622 291952
rect 367730 291864 367910 291952
rect 243214 291648 243394 291736
rect 243502 291648 243682 291736
rect 243790 291648 243970 291736
rect 244078 291648 244258 291736
rect 244366 291648 244546 291736
rect 244654 291648 244834 291736
rect 244942 291648 245122 291736
rect 245230 291648 245410 291736
rect 245664 291648 245844 291736
rect 245952 291648 246132 291736
rect 246240 291648 246420 291736
rect 246528 291648 246708 291736
rect 246816 291648 246996 291736
rect 247104 291648 247284 291736
rect 247392 291648 247572 291736
rect 247680 291648 247860 291736
rect 248114 291648 248294 291736
rect 248402 291648 248582 291736
rect 248690 291648 248870 291736
rect 248978 291648 249158 291736
rect 249266 291648 249446 291736
rect 249554 291648 249734 291736
rect 249842 291648 250022 291736
rect 250130 291648 250310 291736
rect 250564 291648 250744 291736
rect 250852 291648 251032 291736
rect 251140 291648 251320 291736
rect 251428 291648 251608 291736
rect 251716 291648 251896 291736
rect 252004 291648 252184 291736
rect 252292 291648 252472 291736
rect 252580 291648 252760 291736
rect 253014 291648 253194 291736
rect 253302 291648 253482 291736
rect 253590 291648 253770 291736
rect 253878 291648 254058 291736
rect 254166 291648 254346 291736
rect 254454 291648 254634 291736
rect 254742 291648 254922 291736
rect 255030 291648 255210 291736
rect 255464 291648 255644 291736
rect 255752 291648 255932 291736
rect 256040 291648 256220 291736
rect 256328 291648 256508 291736
rect 256616 291648 256796 291736
rect 256904 291648 257084 291736
rect 257192 291648 257372 291736
rect 257480 291648 257660 291736
rect 257914 291648 258094 291736
rect 258202 291648 258382 291736
rect 258490 291648 258670 291736
rect 258778 291648 258958 291736
rect 259066 291648 259246 291736
rect 259354 291648 259534 291736
rect 259642 291648 259822 291736
rect 259930 291648 260110 291736
rect 260364 291648 260544 291736
rect 260652 291648 260832 291736
rect 260940 291648 261120 291736
rect 261228 291648 261408 291736
rect 261516 291648 261696 291736
rect 261804 291648 261984 291736
rect 262092 291648 262272 291736
rect 262380 291648 262560 291736
rect 262814 291648 262994 291736
rect 263102 291648 263282 291736
rect 263390 291648 263570 291736
rect 263678 291648 263858 291736
rect 263966 291648 264146 291736
rect 264254 291648 264434 291736
rect 264542 291648 264722 291736
rect 264830 291648 265010 291736
rect 265264 291648 265444 291736
rect 265552 291648 265732 291736
rect 265840 291648 266020 291736
rect 266128 291648 266308 291736
rect 266416 291648 266596 291736
rect 266704 291648 266884 291736
rect 266992 291648 267172 291736
rect 267280 291648 267460 291736
rect 267714 291648 267894 291736
rect 268002 291648 268182 291736
rect 268290 291648 268470 291736
rect 268578 291648 268758 291736
rect 268866 291648 269046 291736
rect 269154 291648 269334 291736
rect 269442 291648 269622 291736
rect 269730 291648 269910 291736
rect 270164 291648 270344 291736
rect 270452 291648 270632 291736
rect 270740 291648 270920 291736
rect 271028 291648 271208 291736
rect 271316 291648 271496 291736
rect 271604 291648 271784 291736
rect 271892 291648 272072 291736
rect 272180 291648 272360 291736
rect 272614 291648 272794 291736
rect 272902 291648 273082 291736
rect 273190 291648 273370 291736
rect 273478 291648 273658 291736
rect 273766 291648 273946 291736
rect 274054 291648 274234 291736
rect 274342 291648 274522 291736
rect 274630 291648 274810 291736
rect 275064 291648 275244 291736
rect 275352 291648 275532 291736
rect 275640 291648 275820 291736
rect 275928 291648 276108 291736
rect 276216 291648 276396 291736
rect 276504 291648 276684 291736
rect 276792 291648 276972 291736
rect 277080 291648 277260 291736
rect 277514 291648 277694 291736
rect 277802 291648 277982 291736
rect 278090 291648 278270 291736
rect 278378 291648 278558 291736
rect 278666 291648 278846 291736
rect 278954 291648 279134 291736
rect 279242 291648 279422 291736
rect 279530 291648 279710 291736
rect 279964 291648 280144 291736
rect 280252 291648 280432 291736
rect 280540 291648 280720 291736
rect 280828 291648 281008 291736
rect 281116 291648 281296 291736
rect 281404 291648 281584 291736
rect 281692 291648 281872 291736
rect 281980 291648 282160 291736
rect 282414 291648 282594 291736
rect 282702 291648 282882 291736
rect 282990 291648 283170 291736
rect 283278 291648 283458 291736
rect 283566 291648 283746 291736
rect 283854 291648 284034 291736
rect 284142 291648 284322 291736
rect 284430 291648 284610 291736
rect 284864 291648 285044 291736
rect 285152 291648 285332 291736
rect 285440 291648 285620 291736
rect 285728 291648 285908 291736
rect 286016 291648 286196 291736
rect 286304 291648 286484 291736
rect 286592 291648 286772 291736
rect 286880 291648 287060 291736
rect 287314 291648 287494 291736
rect 287602 291648 287782 291736
rect 287890 291648 288070 291736
rect 288178 291648 288358 291736
rect 288466 291648 288646 291736
rect 288754 291648 288934 291736
rect 289042 291648 289222 291736
rect 289330 291648 289510 291736
rect 289764 291648 289944 291736
rect 290052 291648 290232 291736
rect 290340 291648 290520 291736
rect 290628 291648 290808 291736
rect 290916 291648 291096 291736
rect 291204 291648 291384 291736
rect 291492 291648 291672 291736
rect 291780 291648 291960 291736
rect 292214 291648 292394 291736
rect 292502 291648 292682 291736
rect 292790 291648 292970 291736
rect 293078 291648 293258 291736
rect 293366 291648 293546 291736
rect 293654 291648 293834 291736
rect 293942 291648 294122 291736
rect 294230 291648 294410 291736
rect 294664 291648 294844 291736
rect 294952 291648 295132 291736
rect 295240 291648 295420 291736
rect 295528 291648 295708 291736
rect 295816 291648 295996 291736
rect 296104 291648 296284 291736
rect 296392 291648 296572 291736
rect 296680 291648 296860 291736
rect 297114 291648 297294 291736
rect 297402 291648 297582 291736
rect 297690 291648 297870 291736
rect 297978 291648 298158 291736
rect 298266 291648 298446 291736
rect 298554 291648 298734 291736
rect 298842 291648 299022 291736
rect 299130 291648 299310 291736
rect 299564 291648 299744 291736
rect 299852 291648 300032 291736
rect 300140 291648 300320 291736
rect 300428 291648 300608 291736
rect 300716 291648 300896 291736
rect 301004 291648 301184 291736
rect 301292 291648 301472 291736
rect 301580 291648 301760 291736
rect 302014 291648 302194 291736
rect 302302 291648 302482 291736
rect 302590 291648 302770 291736
rect 302878 291648 303058 291736
rect 303166 291648 303346 291736
rect 303454 291648 303634 291736
rect 303742 291648 303922 291736
rect 304030 291648 304210 291736
rect 304464 291648 304644 291736
rect 304752 291648 304932 291736
rect 305040 291648 305220 291736
rect 305328 291648 305508 291736
rect 305616 291648 305796 291736
rect 305904 291648 306084 291736
rect 306192 291648 306372 291736
rect 306480 291648 306660 291736
rect 306914 291648 307094 291736
rect 307202 291648 307382 291736
rect 307490 291648 307670 291736
rect 307778 291648 307958 291736
rect 308066 291648 308246 291736
rect 308354 291648 308534 291736
rect 308642 291648 308822 291736
rect 308930 291648 309110 291736
rect 309364 291648 309544 291736
rect 309652 291648 309832 291736
rect 309940 291648 310120 291736
rect 310228 291648 310408 291736
rect 310516 291648 310696 291736
rect 310804 291648 310984 291736
rect 311092 291648 311272 291736
rect 311380 291648 311560 291736
rect 311814 291648 311994 291736
rect 312102 291648 312282 291736
rect 312390 291648 312570 291736
rect 312678 291648 312858 291736
rect 312966 291648 313146 291736
rect 313254 291648 313434 291736
rect 313542 291648 313722 291736
rect 313830 291648 314010 291736
rect 314264 291648 314444 291736
rect 314552 291648 314732 291736
rect 314840 291648 315020 291736
rect 315128 291648 315308 291736
rect 315416 291648 315596 291736
rect 315704 291648 315884 291736
rect 315992 291648 316172 291736
rect 316280 291648 316460 291736
rect 316714 291648 316894 291736
rect 317002 291648 317182 291736
rect 317290 291648 317470 291736
rect 317578 291648 317758 291736
rect 317866 291648 318046 291736
rect 318154 291648 318334 291736
rect 318442 291648 318622 291736
rect 318730 291648 318910 291736
rect 319164 291648 319344 291736
rect 319452 291648 319632 291736
rect 319740 291648 319920 291736
rect 320028 291648 320208 291736
rect 320316 291648 320496 291736
rect 320604 291648 320784 291736
rect 320892 291648 321072 291736
rect 321180 291648 321360 291736
rect 321614 291648 321794 291736
rect 321902 291648 322082 291736
rect 322190 291648 322370 291736
rect 322478 291648 322658 291736
rect 322766 291648 322946 291736
rect 323054 291648 323234 291736
rect 323342 291648 323522 291736
rect 323630 291648 323810 291736
rect 324064 291648 324244 291736
rect 324352 291648 324532 291736
rect 324640 291648 324820 291736
rect 324928 291648 325108 291736
rect 325216 291648 325396 291736
rect 325504 291648 325684 291736
rect 325792 291648 325972 291736
rect 326080 291648 326260 291736
rect 326514 291648 326694 291736
rect 326802 291648 326982 291736
rect 327090 291648 327270 291736
rect 327378 291648 327558 291736
rect 327666 291648 327846 291736
rect 327954 291648 328134 291736
rect 328242 291648 328422 291736
rect 328530 291648 328710 291736
rect 328964 291648 329144 291736
rect 329252 291648 329432 291736
rect 329540 291648 329720 291736
rect 329828 291648 330008 291736
rect 330116 291648 330296 291736
rect 330404 291648 330584 291736
rect 330692 291648 330872 291736
rect 330980 291648 331160 291736
rect 331414 291648 331594 291736
rect 331702 291648 331882 291736
rect 331990 291648 332170 291736
rect 332278 291648 332458 291736
rect 332566 291648 332746 291736
rect 332854 291648 333034 291736
rect 333142 291648 333322 291736
rect 333430 291648 333610 291736
rect 333864 291648 334044 291736
rect 334152 291648 334332 291736
rect 334440 291648 334620 291736
rect 334728 291648 334908 291736
rect 335016 291648 335196 291736
rect 335304 291648 335484 291736
rect 335592 291648 335772 291736
rect 335880 291648 336060 291736
rect 336314 291648 336494 291736
rect 336602 291648 336782 291736
rect 336890 291648 337070 291736
rect 337178 291648 337358 291736
rect 337466 291648 337646 291736
rect 337754 291648 337934 291736
rect 338042 291648 338222 291736
rect 338330 291648 338510 291736
rect 338764 291648 338944 291736
rect 339052 291648 339232 291736
rect 339340 291648 339520 291736
rect 339628 291648 339808 291736
rect 339916 291648 340096 291736
rect 340204 291648 340384 291736
rect 340492 291648 340672 291736
rect 340780 291648 340960 291736
rect 341214 291648 341394 291736
rect 341502 291648 341682 291736
rect 341790 291648 341970 291736
rect 342078 291648 342258 291736
rect 342366 291648 342546 291736
rect 342654 291648 342834 291736
rect 342942 291648 343122 291736
rect 343230 291648 343410 291736
rect 343664 291648 343844 291736
rect 343952 291648 344132 291736
rect 344240 291648 344420 291736
rect 344528 291648 344708 291736
rect 344816 291648 344996 291736
rect 345104 291648 345284 291736
rect 345392 291648 345572 291736
rect 345680 291648 345860 291736
rect 346114 291648 346294 291736
rect 346402 291648 346582 291736
rect 346690 291648 346870 291736
rect 346978 291648 347158 291736
rect 347266 291648 347446 291736
rect 347554 291648 347734 291736
rect 347842 291648 348022 291736
rect 348130 291648 348310 291736
rect 348564 291648 348744 291736
rect 348852 291648 349032 291736
rect 349140 291648 349320 291736
rect 349428 291648 349608 291736
rect 349716 291648 349896 291736
rect 350004 291648 350184 291736
rect 350292 291648 350472 291736
rect 350580 291648 350760 291736
rect 351014 291648 351194 291736
rect 351302 291648 351482 291736
rect 351590 291648 351770 291736
rect 351878 291648 352058 291736
rect 352166 291648 352346 291736
rect 352454 291648 352634 291736
rect 352742 291648 352922 291736
rect 353030 291648 353210 291736
rect 353464 291648 353644 291736
rect 353752 291648 353932 291736
rect 354040 291648 354220 291736
rect 354328 291648 354508 291736
rect 354616 291648 354796 291736
rect 354904 291648 355084 291736
rect 355192 291648 355372 291736
rect 355480 291648 355660 291736
rect 355914 291648 356094 291736
rect 356202 291648 356382 291736
rect 356490 291648 356670 291736
rect 356778 291648 356958 291736
rect 357066 291648 357246 291736
rect 357354 291648 357534 291736
rect 357642 291648 357822 291736
rect 357930 291648 358110 291736
rect 358364 291648 358544 291736
rect 358652 291648 358832 291736
rect 358940 291648 359120 291736
rect 359228 291648 359408 291736
rect 359516 291648 359696 291736
rect 359804 291648 359984 291736
rect 360092 291648 360272 291736
rect 360380 291648 360560 291736
rect 360814 291648 360994 291736
rect 361102 291648 361282 291736
rect 361390 291648 361570 291736
rect 361678 291648 361858 291736
rect 361966 291648 362146 291736
rect 362254 291648 362434 291736
rect 362542 291648 362722 291736
rect 362830 291648 363010 291736
rect 363264 291648 363444 291736
rect 363552 291648 363732 291736
rect 363840 291648 364020 291736
rect 364128 291648 364308 291736
rect 364416 291648 364596 291736
rect 364704 291648 364884 291736
rect 364992 291648 365172 291736
rect 365280 291648 365460 291736
rect 365714 291648 365894 291736
rect 366002 291648 366182 291736
rect 366290 291648 366470 291736
rect 366578 291648 366758 291736
rect 366866 291648 367046 291736
rect 367154 291648 367334 291736
rect 367442 291648 367622 291736
rect 367730 291648 367910 291736
rect 243214 291172 243394 291260
rect 243502 291172 243682 291260
rect 243790 291172 243970 291260
rect 244078 291172 244258 291260
rect 244366 291172 244546 291260
rect 244654 291172 244834 291260
rect 244942 291172 245122 291260
rect 245230 291172 245410 291260
rect 245664 291172 245844 291260
rect 245952 291172 246132 291260
rect 246240 291172 246420 291260
rect 246528 291172 246708 291260
rect 246816 291172 246996 291260
rect 247104 291172 247284 291260
rect 247392 291172 247572 291260
rect 247680 291172 247860 291260
rect 248114 291172 248294 291260
rect 248402 291172 248582 291260
rect 248690 291172 248870 291260
rect 248978 291172 249158 291260
rect 249266 291172 249446 291260
rect 249554 291172 249734 291260
rect 249842 291172 250022 291260
rect 250130 291172 250310 291260
rect 250564 291172 250744 291260
rect 250852 291172 251032 291260
rect 251140 291172 251320 291260
rect 251428 291172 251608 291260
rect 251716 291172 251896 291260
rect 252004 291172 252184 291260
rect 252292 291172 252472 291260
rect 252580 291172 252760 291260
rect 253014 291172 253194 291260
rect 253302 291172 253482 291260
rect 253590 291172 253770 291260
rect 253878 291172 254058 291260
rect 254166 291172 254346 291260
rect 254454 291172 254634 291260
rect 254742 291172 254922 291260
rect 255030 291172 255210 291260
rect 255464 291172 255644 291260
rect 255752 291172 255932 291260
rect 256040 291172 256220 291260
rect 256328 291172 256508 291260
rect 256616 291172 256796 291260
rect 256904 291172 257084 291260
rect 257192 291172 257372 291260
rect 257480 291172 257660 291260
rect 257914 291172 258094 291260
rect 258202 291172 258382 291260
rect 258490 291172 258670 291260
rect 258778 291172 258958 291260
rect 259066 291172 259246 291260
rect 259354 291172 259534 291260
rect 259642 291172 259822 291260
rect 259930 291172 260110 291260
rect 260364 291172 260544 291260
rect 260652 291172 260832 291260
rect 260940 291172 261120 291260
rect 261228 291172 261408 291260
rect 261516 291172 261696 291260
rect 261804 291172 261984 291260
rect 262092 291172 262272 291260
rect 262380 291172 262560 291260
rect 262814 291172 262994 291260
rect 263102 291172 263282 291260
rect 263390 291172 263570 291260
rect 263678 291172 263858 291260
rect 263966 291172 264146 291260
rect 264254 291172 264434 291260
rect 264542 291172 264722 291260
rect 264830 291172 265010 291260
rect 265264 291172 265444 291260
rect 265552 291172 265732 291260
rect 265840 291172 266020 291260
rect 266128 291172 266308 291260
rect 266416 291172 266596 291260
rect 266704 291172 266884 291260
rect 266992 291172 267172 291260
rect 267280 291172 267460 291260
rect 267714 291172 267894 291260
rect 268002 291172 268182 291260
rect 268290 291172 268470 291260
rect 268578 291172 268758 291260
rect 268866 291172 269046 291260
rect 269154 291172 269334 291260
rect 269442 291172 269622 291260
rect 269730 291172 269910 291260
rect 270164 291172 270344 291260
rect 270452 291172 270632 291260
rect 270740 291172 270920 291260
rect 271028 291172 271208 291260
rect 271316 291172 271496 291260
rect 271604 291172 271784 291260
rect 271892 291172 272072 291260
rect 272180 291172 272360 291260
rect 272614 291172 272794 291260
rect 272902 291172 273082 291260
rect 273190 291172 273370 291260
rect 273478 291172 273658 291260
rect 273766 291172 273946 291260
rect 274054 291172 274234 291260
rect 274342 291172 274522 291260
rect 274630 291172 274810 291260
rect 275064 291172 275244 291260
rect 275352 291172 275532 291260
rect 275640 291172 275820 291260
rect 275928 291172 276108 291260
rect 276216 291172 276396 291260
rect 276504 291172 276684 291260
rect 276792 291172 276972 291260
rect 277080 291172 277260 291260
rect 277514 291172 277694 291260
rect 277802 291172 277982 291260
rect 278090 291172 278270 291260
rect 278378 291172 278558 291260
rect 278666 291172 278846 291260
rect 278954 291172 279134 291260
rect 279242 291172 279422 291260
rect 279530 291172 279710 291260
rect 279964 291172 280144 291260
rect 280252 291172 280432 291260
rect 280540 291172 280720 291260
rect 280828 291172 281008 291260
rect 281116 291172 281296 291260
rect 281404 291172 281584 291260
rect 281692 291172 281872 291260
rect 281980 291172 282160 291260
rect 282414 291172 282594 291260
rect 282702 291172 282882 291260
rect 282990 291172 283170 291260
rect 283278 291172 283458 291260
rect 283566 291172 283746 291260
rect 283854 291172 284034 291260
rect 284142 291172 284322 291260
rect 284430 291172 284610 291260
rect 284864 291172 285044 291260
rect 285152 291172 285332 291260
rect 285440 291172 285620 291260
rect 285728 291172 285908 291260
rect 286016 291172 286196 291260
rect 286304 291172 286484 291260
rect 286592 291172 286772 291260
rect 286880 291172 287060 291260
rect 287314 291172 287494 291260
rect 287602 291172 287782 291260
rect 287890 291172 288070 291260
rect 288178 291172 288358 291260
rect 288466 291172 288646 291260
rect 288754 291172 288934 291260
rect 289042 291172 289222 291260
rect 289330 291172 289510 291260
rect 289764 291172 289944 291260
rect 290052 291172 290232 291260
rect 290340 291172 290520 291260
rect 290628 291172 290808 291260
rect 290916 291172 291096 291260
rect 291204 291172 291384 291260
rect 291492 291172 291672 291260
rect 291780 291172 291960 291260
rect 292214 291172 292394 291260
rect 292502 291172 292682 291260
rect 292790 291172 292970 291260
rect 293078 291172 293258 291260
rect 293366 291172 293546 291260
rect 293654 291172 293834 291260
rect 293942 291172 294122 291260
rect 294230 291172 294410 291260
rect 294664 291172 294844 291260
rect 294952 291172 295132 291260
rect 295240 291172 295420 291260
rect 295528 291172 295708 291260
rect 295816 291172 295996 291260
rect 296104 291172 296284 291260
rect 296392 291172 296572 291260
rect 296680 291172 296860 291260
rect 297114 291172 297294 291260
rect 297402 291172 297582 291260
rect 297690 291172 297870 291260
rect 297978 291172 298158 291260
rect 298266 291172 298446 291260
rect 298554 291172 298734 291260
rect 298842 291172 299022 291260
rect 299130 291172 299310 291260
rect 299564 291172 299744 291260
rect 299852 291172 300032 291260
rect 300140 291172 300320 291260
rect 300428 291172 300608 291260
rect 300716 291172 300896 291260
rect 301004 291172 301184 291260
rect 301292 291172 301472 291260
rect 301580 291172 301760 291260
rect 302014 291172 302194 291260
rect 302302 291172 302482 291260
rect 302590 291172 302770 291260
rect 302878 291172 303058 291260
rect 303166 291172 303346 291260
rect 303454 291172 303634 291260
rect 303742 291172 303922 291260
rect 304030 291172 304210 291260
rect 304464 291172 304644 291260
rect 304752 291172 304932 291260
rect 305040 291172 305220 291260
rect 305328 291172 305508 291260
rect 305616 291172 305796 291260
rect 305904 291172 306084 291260
rect 306192 291172 306372 291260
rect 306480 291172 306660 291260
rect 306914 291172 307094 291260
rect 307202 291172 307382 291260
rect 307490 291172 307670 291260
rect 307778 291172 307958 291260
rect 308066 291172 308246 291260
rect 308354 291172 308534 291260
rect 308642 291172 308822 291260
rect 308930 291172 309110 291260
rect 309364 291172 309544 291260
rect 309652 291172 309832 291260
rect 309940 291172 310120 291260
rect 310228 291172 310408 291260
rect 310516 291172 310696 291260
rect 310804 291172 310984 291260
rect 311092 291172 311272 291260
rect 311380 291172 311560 291260
rect 311814 291172 311994 291260
rect 312102 291172 312282 291260
rect 312390 291172 312570 291260
rect 312678 291172 312858 291260
rect 312966 291172 313146 291260
rect 313254 291172 313434 291260
rect 313542 291172 313722 291260
rect 313830 291172 314010 291260
rect 314264 291172 314444 291260
rect 314552 291172 314732 291260
rect 314840 291172 315020 291260
rect 315128 291172 315308 291260
rect 315416 291172 315596 291260
rect 315704 291172 315884 291260
rect 315992 291172 316172 291260
rect 316280 291172 316460 291260
rect 316714 291172 316894 291260
rect 317002 291172 317182 291260
rect 317290 291172 317470 291260
rect 317578 291172 317758 291260
rect 317866 291172 318046 291260
rect 318154 291172 318334 291260
rect 318442 291172 318622 291260
rect 318730 291172 318910 291260
rect 319164 291172 319344 291260
rect 319452 291172 319632 291260
rect 319740 291172 319920 291260
rect 320028 291172 320208 291260
rect 320316 291172 320496 291260
rect 320604 291172 320784 291260
rect 320892 291172 321072 291260
rect 321180 291172 321360 291260
rect 321614 291172 321794 291260
rect 321902 291172 322082 291260
rect 322190 291172 322370 291260
rect 322478 291172 322658 291260
rect 322766 291172 322946 291260
rect 323054 291172 323234 291260
rect 323342 291172 323522 291260
rect 323630 291172 323810 291260
rect 324064 291172 324244 291260
rect 324352 291172 324532 291260
rect 324640 291172 324820 291260
rect 324928 291172 325108 291260
rect 325216 291172 325396 291260
rect 325504 291172 325684 291260
rect 325792 291172 325972 291260
rect 326080 291172 326260 291260
rect 326514 291172 326694 291260
rect 326802 291172 326982 291260
rect 327090 291172 327270 291260
rect 327378 291172 327558 291260
rect 327666 291172 327846 291260
rect 327954 291172 328134 291260
rect 328242 291172 328422 291260
rect 328530 291172 328710 291260
rect 328964 291172 329144 291260
rect 329252 291172 329432 291260
rect 329540 291172 329720 291260
rect 329828 291172 330008 291260
rect 330116 291172 330296 291260
rect 330404 291172 330584 291260
rect 330692 291172 330872 291260
rect 330980 291172 331160 291260
rect 331414 291172 331594 291260
rect 331702 291172 331882 291260
rect 331990 291172 332170 291260
rect 332278 291172 332458 291260
rect 332566 291172 332746 291260
rect 332854 291172 333034 291260
rect 333142 291172 333322 291260
rect 333430 291172 333610 291260
rect 333864 291172 334044 291260
rect 334152 291172 334332 291260
rect 334440 291172 334620 291260
rect 334728 291172 334908 291260
rect 335016 291172 335196 291260
rect 335304 291172 335484 291260
rect 335592 291172 335772 291260
rect 335880 291172 336060 291260
rect 336314 291172 336494 291260
rect 336602 291172 336782 291260
rect 336890 291172 337070 291260
rect 337178 291172 337358 291260
rect 337466 291172 337646 291260
rect 337754 291172 337934 291260
rect 338042 291172 338222 291260
rect 338330 291172 338510 291260
rect 338764 291172 338944 291260
rect 339052 291172 339232 291260
rect 339340 291172 339520 291260
rect 339628 291172 339808 291260
rect 339916 291172 340096 291260
rect 340204 291172 340384 291260
rect 340492 291172 340672 291260
rect 340780 291172 340960 291260
rect 341214 291172 341394 291260
rect 341502 291172 341682 291260
rect 341790 291172 341970 291260
rect 342078 291172 342258 291260
rect 342366 291172 342546 291260
rect 342654 291172 342834 291260
rect 342942 291172 343122 291260
rect 343230 291172 343410 291260
rect 343664 291172 343844 291260
rect 343952 291172 344132 291260
rect 344240 291172 344420 291260
rect 344528 291172 344708 291260
rect 344816 291172 344996 291260
rect 345104 291172 345284 291260
rect 345392 291172 345572 291260
rect 345680 291172 345860 291260
rect 346114 291172 346294 291260
rect 346402 291172 346582 291260
rect 346690 291172 346870 291260
rect 346978 291172 347158 291260
rect 347266 291172 347446 291260
rect 347554 291172 347734 291260
rect 347842 291172 348022 291260
rect 348130 291172 348310 291260
rect 348564 291172 348744 291260
rect 348852 291172 349032 291260
rect 349140 291172 349320 291260
rect 349428 291172 349608 291260
rect 349716 291172 349896 291260
rect 350004 291172 350184 291260
rect 350292 291172 350472 291260
rect 350580 291172 350760 291260
rect 351014 291172 351194 291260
rect 351302 291172 351482 291260
rect 351590 291172 351770 291260
rect 351878 291172 352058 291260
rect 352166 291172 352346 291260
rect 352454 291172 352634 291260
rect 352742 291172 352922 291260
rect 353030 291172 353210 291260
rect 353464 291172 353644 291260
rect 353752 291172 353932 291260
rect 354040 291172 354220 291260
rect 354328 291172 354508 291260
rect 354616 291172 354796 291260
rect 354904 291172 355084 291260
rect 355192 291172 355372 291260
rect 355480 291172 355660 291260
rect 355914 291172 356094 291260
rect 356202 291172 356382 291260
rect 356490 291172 356670 291260
rect 356778 291172 356958 291260
rect 357066 291172 357246 291260
rect 357354 291172 357534 291260
rect 357642 291172 357822 291260
rect 357930 291172 358110 291260
rect 358364 291172 358544 291260
rect 358652 291172 358832 291260
rect 358940 291172 359120 291260
rect 359228 291172 359408 291260
rect 359516 291172 359696 291260
rect 359804 291172 359984 291260
rect 360092 291172 360272 291260
rect 360380 291172 360560 291260
rect 360814 291172 360994 291260
rect 361102 291172 361282 291260
rect 361390 291172 361570 291260
rect 361678 291172 361858 291260
rect 361966 291172 362146 291260
rect 362254 291172 362434 291260
rect 362542 291172 362722 291260
rect 362830 291172 363010 291260
rect 363264 291172 363444 291260
rect 363552 291172 363732 291260
rect 363840 291172 364020 291260
rect 364128 291172 364308 291260
rect 364416 291172 364596 291260
rect 364704 291172 364884 291260
rect 364992 291172 365172 291260
rect 365280 291172 365460 291260
rect 365714 291172 365894 291260
rect 366002 291172 366182 291260
rect 366290 291172 366470 291260
rect 366578 291172 366758 291260
rect 366866 291172 367046 291260
rect 367154 291172 367334 291260
rect 367442 291172 367622 291260
rect 367730 291172 367910 291260
rect 243214 290698 243394 290786
rect 243502 290698 243682 290786
rect 243790 290698 243970 290786
rect 244078 290698 244258 290786
rect 244366 290698 244546 290786
rect 244654 290698 244834 290786
rect 244942 290698 245122 290786
rect 245230 290698 245410 290786
rect 245664 290698 245844 290786
rect 245952 290698 246132 290786
rect 246240 290698 246420 290786
rect 246528 290698 246708 290786
rect 246816 290698 246996 290786
rect 247104 290698 247284 290786
rect 247392 290698 247572 290786
rect 247680 290698 247860 290786
rect 248114 290698 248294 290786
rect 248402 290698 248582 290786
rect 248690 290698 248870 290786
rect 248978 290698 249158 290786
rect 249266 290698 249446 290786
rect 249554 290698 249734 290786
rect 249842 290698 250022 290786
rect 250130 290698 250310 290786
rect 250564 290698 250744 290786
rect 250852 290698 251032 290786
rect 251140 290698 251320 290786
rect 251428 290698 251608 290786
rect 251716 290698 251896 290786
rect 252004 290698 252184 290786
rect 252292 290698 252472 290786
rect 252580 290698 252760 290786
rect 253014 290698 253194 290786
rect 253302 290698 253482 290786
rect 253590 290698 253770 290786
rect 253878 290698 254058 290786
rect 254166 290698 254346 290786
rect 254454 290698 254634 290786
rect 254742 290698 254922 290786
rect 255030 290698 255210 290786
rect 255464 290698 255644 290786
rect 255752 290698 255932 290786
rect 256040 290698 256220 290786
rect 256328 290698 256508 290786
rect 256616 290698 256796 290786
rect 256904 290698 257084 290786
rect 257192 290698 257372 290786
rect 257480 290698 257660 290786
rect 257914 290698 258094 290786
rect 258202 290698 258382 290786
rect 258490 290698 258670 290786
rect 258778 290698 258958 290786
rect 259066 290698 259246 290786
rect 259354 290698 259534 290786
rect 259642 290698 259822 290786
rect 259930 290698 260110 290786
rect 260364 290698 260544 290786
rect 260652 290698 260832 290786
rect 260940 290698 261120 290786
rect 261228 290698 261408 290786
rect 261516 290698 261696 290786
rect 261804 290698 261984 290786
rect 262092 290698 262272 290786
rect 262380 290698 262560 290786
rect 262814 290698 262994 290786
rect 263102 290698 263282 290786
rect 263390 290698 263570 290786
rect 263678 290698 263858 290786
rect 263966 290698 264146 290786
rect 264254 290698 264434 290786
rect 264542 290698 264722 290786
rect 264830 290698 265010 290786
rect 265264 290698 265444 290786
rect 265552 290698 265732 290786
rect 265840 290698 266020 290786
rect 266128 290698 266308 290786
rect 266416 290698 266596 290786
rect 266704 290698 266884 290786
rect 266992 290698 267172 290786
rect 267280 290698 267460 290786
rect 267714 290698 267894 290786
rect 268002 290698 268182 290786
rect 268290 290698 268470 290786
rect 268578 290698 268758 290786
rect 268866 290698 269046 290786
rect 269154 290698 269334 290786
rect 269442 290698 269622 290786
rect 269730 290698 269910 290786
rect 270164 290698 270344 290786
rect 270452 290698 270632 290786
rect 270740 290698 270920 290786
rect 271028 290698 271208 290786
rect 271316 290698 271496 290786
rect 271604 290698 271784 290786
rect 271892 290698 272072 290786
rect 272180 290698 272360 290786
rect 272614 290698 272794 290786
rect 272902 290698 273082 290786
rect 273190 290698 273370 290786
rect 273478 290698 273658 290786
rect 273766 290698 273946 290786
rect 274054 290698 274234 290786
rect 274342 290698 274522 290786
rect 274630 290698 274810 290786
rect 275064 290698 275244 290786
rect 275352 290698 275532 290786
rect 275640 290698 275820 290786
rect 275928 290698 276108 290786
rect 276216 290698 276396 290786
rect 276504 290698 276684 290786
rect 276792 290698 276972 290786
rect 277080 290698 277260 290786
rect 277514 290698 277694 290786
rect 277802 290698 277982 290786
rect 278090 290698 278270 290786
rect 278378 290698 278558 290786
rect 278666 290698 278846 290786
rect 278954 290698 279134 290786
rect 279242 290698 279422 290786
rect 279530 290698 279710 290786
rect 279964 290698 280144 290786
rect 280252 290698 280432 290786
rect 280540 290698 280720 290786
rect 280828 290698 281008 290786
rect 281116 290698 281296 290786
rect 281404 290698 281584 290786
rect 281692 290698 281872 290786
rect 281980 290698 282160 290786
rect 282414 290698 282594 290786
rect 282702 290698 282882 290786
rect 282990 290698 283170 290786
rect 283278 290698 283458 290786
rect 283566 290698 283746 290786
rect 283854 290698 284034 290786
rect 284142 290698 284322 290786
rect 284430 290698 284610 290786
rect 284864 290698 285044 290786
rect 285152 290698 285332 290786
rect 285440 290698 285620 290786
rect 285728 290698 285908 290786
rect 286016 290698 286196 290786
rect 286304 290698 286484 290786
rect 286592 290698 286772 290786
rect 286880 290698 287060 290786
rect 287314 290698 287494 290786
rect 287602 290698 287782 290786
rect 287890 290698 288070 290786
rect 288178 290698 288358 290786
rect 288466 290698 288646 290786
rect 288754 290698 288934 290786
rect 289042 290698 289222 290786
rect 289330 290698 289510 290786
rect 289764 290698 289944 290786
rect 290052 290698 290232 290786
rect 290340 290698 290520 290786
rect 290628 290698 290808 290786
rect 290916 290698 291096 290786
rect 291204 290698 291384 290786
rect 291492 290698 291672 290786
rect 291780 290698 291960 290786
rect 292214 290698 292394 290786
rect 292502 290698 292682 290786
rect 292790 290698 292970 290786
rect 293078 290698 293258 290786
rect 293366 290698 293546 290786
rect 293654 290698 293834 290786
rect 293942 290698 294122 290786
rect 294230 290698 294410 290786
rect 294664 290698 294844 290786
rect 294952 290698 295132 290786
rect 295240 290698 295420 290786
rect 295528 290698 295708 290786
rect 295816 290698 295996 290786
rect 296104 290698 296284 290786
rect 296392 290698 296572 290786
rect 296680 290698 296860 290786
rect 297114 290698 297294 290786
rect 297402 290698 297582 290786
rect 297690 290698 297870 290786
rect 297978 290698 298158 290786
rect 298266 290698 298446 290786
rect 298554 290698 298734 290786
rect 298842 290698 299022 290786
rect 299130 290698 299310 290786
rect 299564 290698 299744 290786
rect 299852 290698 300032 290786
rect 300140 290698 300320 290786
rect 300428 290698 300608 290786
rect 300716 290698 300896 290786
rect 301004 290698 301184 290786
rect 301292 290698 301472 290786
rect 301580 290698 301760 290786
rect 302014 290698 302194 290786
rect 302302 290698 302482 290786
rect 302590 290698 302770 290786
rect 302878 290698 303058 290786
rect 303166 290698 303346 290786
rect 303454 290698 303634 290786
rect 303742 290698 303922 290786
rect 304030 290698 304210 290786
rect 304464 290698 304644 290786
rect 304752 290698 304932 290786
rect 305040 290698 305220 290786
rect 305328 290698 305508 290786
rect 305616 290698 305796 290786
rect 305904 290698 306084 290786
rect 306192 290698 306372 290786
rect 306480 290698 306660 290786
rect 306914 290698 307094 290786
rect 307202 290698 307382 290786
rect 307490 290698 307670 290786
rect 307778 290698 307958 290786
rect 308066 290698 308246 290786
rect 308354 290698 308534 290786
rect 308642 290698 308822 290786
rect 308930 290698 309110 290786
rect 309364 290698 309544 290786
rect 309652 290698 309832 290786
rect 309940 290698 310120 290786
rect 310228 290698 310408 290786
rect 310516 290698 310696 290786
rect 310804 290698 310984 290786
rect 311092 290698 311272 290786
rect 311380 290698 311560 290786
rect 311814 290698 311994 290786
rect 312102 290698 312282 290786
rect 312390 290698 312570 290786
rect 312678 290698 312858 290786
rect 312966 290698 313146 290786
rect 313254 290698 313434 290786
rect 313542 290698 313722 290786
rect 313830 290698 314010 290786
rect 314264 290698 314444 290786
rect 314552 290698 314732 290786
rect 314840 290698 315020 290786
rect 315128 290698 315308 290786
rect 315416 290698 315596 290786
rect 315704 290698 315884 290786
rect 315992 290698 316172 290786
rect 316280 290698 316460 290786
rect 316714 290698 316894 290786
rect 317002 290698 317182 290786
rect 317290 290698 317470 290786
rect 317578 290698 317758 290786
rect 317866 290698 318046 290786
rect 318154 290698 318334 290786
rect 318442 290698 318622 290786
rect 318730 290698 318910 290786
rect 319164 290698 319344 290786
rect 319452 290698 319632 290786
rect 319740 290698 319920 290786
rect 320028 290698 320208 290786
rect 320316 290698 320496 290786
rect 320604 290698 320784 290786
rect 320892 290698 321072 290786
rect 321180 290698 321360 290786
rect 321614 290698 321794 290786
rect 321902 290698 322082 290786
rect 322190 290698 322370 290786
rect 322478 290698 322658 290786
rect 322766 290698 322946 290786
rect 323054 290698 323234 290786
rect 323342 290698 323522 290786
rect 323630 290698 323810 290786
rect 324064 290698 324244 290786
rect 324352 290698 324532 290786
rect 324640 290698 324820 290786
rect 324928 290698 325108 290786
rect 325216 290698 325396 290786
rect 325504 290698 325684 290786
rect 325792 290698 325972 290786
rect 326080 290698 326260 290786
rect 326514 290698 326694 290786
rect 326802 290698 326982 290786
rect 327090 290698 327270 290786
rect 327378 290698 327558 290786
rect 327666 290698 327846 290786
rect 327954 290698 328134 290786
rect 328242 290698 328422 290786
rect 328530 290698 328710 290786
rect 328964 290698 329144 290786
rect 329252 290698 329432 290786
rect 329540 290698 329720 290786
rect 329828 290698 330008 290786
rect 330116 290698 330296 290786
rect 330404 290698 330584 290786
rect 330692 290698 330872 290786
rect 330980 290698 331160 290786
rect 331414 290698 331594 290786
rect 331702 290698 331882 290786
rect 331990 290698 332170 290786
rect 332278 290698 332458 290786
rect 332566 290698 332746 290786
rect 332854 290698 333034 290786
rect 333142 290698 333322 290786
rect 333430 290698 333610 290786
rect 333864 290698 334044 290786
rect 334152 290698 334332 290786
rect 334440 290698 334620 290786
rect 334728 290698 334908 290786
rect 335016 290698 335196 290786
rect 335304 290698 335484 290786
rect 335592 290698 335772 290786
rect 335880 290698 336060 290786
rect 336314 290698 336494 290786
rect 336602 290698 336782 290786
rect 336890 290698 337070 290786
rect 337178 290698 337358 290786
rect 337466 290698 337646 290786
rect 337754 290698 337934 290786
rect 338042 290698 338222 290786
rect 338330 290698 338510 290786
rect 338764 290698 338944 290786
rect 339052 290698 339232 290786
rect 339340 290698 339520 290786
rect 339628 290698 339808 290786
rect 339916 290698 340096 290786
rect 340204 290698 340384 290786
rect 340492 290698 340672 290786
rect 340780 290698 340960 290786
rect 341214 290698 341394 290786
rect 341502 290698 341682 290786
rect 341790 290698 341970 290786
rect 342078 290698 342258 290786
rect 342366 290698 342546 290786
rect 342654 290698 342834 290786
rect 342942 290698 343122 290786
rect 343230 290698 343410 290786
rect 343664 290698 343844 290786
rect 343952 290698 344132 290786
rect 344240 290698 344420 290786
rect 344528 290698 344708 290786
rect 344816 290698 344996 290786
rect 345104 290698 345284 290786
rect 345392 290698 345572 290786
rect 345680 290698 345860 290786
rect 346114 290698 346294 290786
rect 346402 290698 346582 290786
rect 346690 290698 346870 290786
rect 346978 290698 347158 290786
rect 347266 290698 347446 290786
rect 347554 290698 347734 290786
rect 347842 290698 348022 290786
rect 348130 290698 348310 290786
rect 348564 290698 348744 290786
rect 348852 290698 349032 290786
rect 349140 290698 349320 290786
rect 349428 290698 349608 290786
rect 349716 290698 349896 290786
rect 350004 290698 350184 290786
rect 350292 290698 350472 290786
rect 350580 290698 350760 290786
rect 351014 290698 351194 290786
rect 351302 290698 351482 290786
rect 351590 290698 351770 290786
rect 351878 290698 352058 290786
rect 352166 290698 352346 290786
rect 352454 290698 352634 290786
rect 352742 290698 352922 290786
rect 353030 290698 353210 290786
rect 353464 290698 353644 290786
rect 353752 290698 353932 290786
rect 354040 290698 354220 290786
rect 354328 290698 354508 290786
rect 354616 290698 354796 290786
rect 354904 290698 355084 290786
rect 355192 290698 355372 290786
rect 355480 290698 355660 290786
rect 355914 290698 356094 290786
rect 356202 290698 356382 290786
rect 356490 290698 356670 290786
rect 356778 290698 356958 290786
rect 357066 290698 357246 290786
rect 357354 290698 357534 290786
rect 357642 290698 357822 290786
rect 357930 290698 358110 290786
rect 358364 290698 358544 290786
rect 358652 290698 358832 290786
rect 358940 290698 359120 290786
rect 359228 290698 359408 290786
rect 359516 290698 359696 290786
rect 359804 290698 359984 290786
rect 360092 290698 360272 290786
rect 360380 290698 360560 290786
rect 360814 290698 360994 290786
rect 361102 290698 361282 290786
rect 361390 290698 361570 290786
rect 361678 290698 361858 290786
rect 361966 290698 362146 290786
rect 362254 290698 362434 290786
rect 362542 290698 362722 290786
rect 362830 290698 363010 290786
rect 363264 290698 363444 290786
rect 363552 290698 363732 290786
rect 363840 290698 364020 290786
rect 364128 290698 364308 290786
rect 364416 290698 364596 290786
rect 364704 290698 364884 290786
rect 364992 290698 365172 290786
rect 365280 290698 365460 290786
rect 365714 290698 365894 290786
rect 366002 290698 366182 290786
rect 366290 290698 366470 290786
rect 366578 290698 366758 290786
rect 366866 290698 367046 290786
rect 367154 290698 367334 290786
rect 367442 290698 367622 290786
rect 367730 290698 367910 290786
rect 243214 290222 243394 290310
rect 243502 290222 243682 290310
rect 243790 290222 243970 290310
rect 244078 290222 244258 290310
rect 244366 290222 244546 290310
rect 244654 290222 244834 290310
rect 244942 290222 245122 290310
rect 245230 290222 245410 290310
rect 245664 290222 245844 290310
rect 245952 290222 246132 290310
rect 246240 290222 246420 290310
rect 246528 290222 246708 290310
rect 246816 290222 246996 290310
rect 247104 290222 247284 290310
rect 247392 290222 247572 290310
rect 247680 290222 247860 290310
rect 248114 290222 248294 290310
rect 248402 290222 248582 290310
rect 248690 290222 248870 290310
rect 248978 290222 249158 290310
rect 249266 290222 249446 290310
rect 249554 290222 249734 290310
rect 249842 290222 250022 290310
rect 250130 290222 250310 290310
rect 250564 290222 250744 290310
rect 250852 290222 251032 290310
rect 251140 290222 251320 290310
rect 251428 290222 251608 290310
rect 251716 290222 251896 290310
rect 252004 290222 252184 290310
rect 252292 290222 252472 290310
rect 252580 290222 252760 290310
rect 253014 290222 253194 290310
rect 253302 290222 253482 290310
rect 253590 290222 253770 290310
rect 253878 290222 254058 290310
rect 254166 290222 254346 290310
rect 254454 290222 254634 290310
rect 254742 290222 254922 290310
rect 255030 290222 255210 290310
rect 255464 290222 255644 290310
rect 255752 290222 255932 290310
rect 256040 290222 256220 290310
rect 256328 290222 256508 290310
rect 256616 290222 256796 290310
rect 256904 290222 257084 290310
rect 257192 290222 257372 290310
rect 257480 290222 257660 290310
rect 257914 290222 258094 290310
rect 258202 290222 258382 290310
rect 258490 290222 258670 290310
rect 258778 290222 258958 290310
rect 259066 290222 259246 290310
rect 259354 290222 259534 290310
rect 259642 290222 259822 290310
rect 259930 290222 260110 290310
rect 260364 290222 260544 290310
rect 260652 290222 260832 290310
rect 260940 290222 261120 290310
rect 261228 290222 261408 290310
rect 261516 290222 261696 290310
rect 261804 290222 261984 290310
rect 262092 290222 262272 290310
rect 262380 290222 262560 290310
rect 262814 290222 262994 290310
rect 263102 290222 263282 290310
rect 263390 290222 263570 290310
rect 263678 290222 263858 290310
rect 263966 290222 264146 290310
rect 264254 290222 264434 290310
rect 264542 290222 264722 290310
rect 264830 290222 265010 290310
rect 265264 290222 265444 290310
rect 265552 290222 265732 290310
rect 265840 290222 266020 290310
rect 266128 290222 266308 290310
rect 266416 290222 266596 290310
rect 266704 290222 266884 290310
rect 266992 290222 267172 290310
rect 267280 290222 267460 290310
rect 267714 290222 267894 290310
rect 268002 290222 268182 290310
rect 268290 290222 268470 290310
rect 268578 290222 268758 290310
rect 268866 290222 269046 290310
rect 269154 290222 269334 290310
rect 269442 290222 269622 290310
rect 269730 290222 269910 290310
rect 270164 290222 270344 290310
rect 270452 290222 270632 290310
rect 270740 290222 270920 290310
rect 271028 290222 271208 290310
rect 271316 290222 271496 290310
rect 271604 290222 271784 290310
rect 271892 290222 272072 290310
rect 272180 290222 272360 290310
rect 272614 290222 272794 290310
rect 272902 290222 273082 290310
rect 273190 290222 273370 290310
rect 273478 290222 273658 290310
rect 273766 290222 273946 290310
rect 274054 290222 274234 290310
rect 274342 290222 274522 290310
rect 274630 290222 274810 290310
rect 275064 290222 275244 290310
rect 275352 290222 275532 290310
rect 275640 290222 275820 290310
rect 275928 290222 276108 290310
rect 276216 290222 276396 290310
rect 276504 290222 276684 290310
rect 276792 290222 276972 290310
rect 277080 290222 277260 290310
rect 277514 290222 277694 290310
rect 277802 290222 277982 290310
rect 278090 290222 278270 290310
rect 278378 290222 278558 290310
rect 278666 290222 278846 290310
rect 278954 290222 279134 290310
rect 279242 290222 279422 290310
rect 279530 290222 279710 290310
rect 279964 290222 280144 290310
rect 280252 290222 280432 290310
rect 280540 290222 280720 290310
rect 280828 290222 281008 290310
rect 281116 290222 281296 290310
rect 281404 290222 281584 290310
rect 281692 290222 281872 290310
rect 281980 290222 282160 290310
rect 282414 290222 282594 290310
rect 282702 290222 282882 290310
rect 282990 290222 283170 290310
rect 283278 290222 283458 290310
rect 283566 290222 283746 290310
rect 283854 290222 284034 290310
rect 284142 290222 284322 290310
rect 284430 290222 284610 290310
rect 284864 290222 285044 290310
rect 285152 290222 285332 290310
rect 285440 290222 285620 290310
rect 285728 290222 285908 290310
rect 286016 290222 286196 290310
rect 286304 290222 286484 290310
rect 286592 290222 286772 290310
rect 286880 290222 287060 290310
rect 287314 290222 287494 290310
rect 287602 290222 287782 290310
rect 287890 290222 288070 290310
rect 288178 290222 288358 290310
rect 288466 290222 288646 290310
rect 288754 290222 288934 290310
rect 289042 290222 289222 290310
rect 289330 290222 289510 290310
rect 289764 290222 289944 290310
rect 290052 290222 290232 290310
rect 290340 290222 290520 290310
rect 290628 290222 290808 290310
rect 290916 290222 291096 290310
rect 291204 290222 291384 290310
rect 291492 290222 291672 290310
rect 291780 290222 291960 290310
rect 292214 290222 292394 290310
rect 292502 290222 292682 290310
rect 292790 290222 292970 290310
rect 293078 290222 293258 290310
rect 293366 290222 293546 290310
rect 293654 290222 293834 290310
rect 293942 290222 294122 290310
rect 294230 290222 294410 290310
rect 294664 290222 294844 290310
rect 294952 290222 295132 290310
rect 295240 290222 295420 290310
rect 295528 290222 295708 290310
rect 295816 290222 295996 290310
rect 296104 290222 296284 290310
rect 296392 290222 296572 290310
rect 296680 290222 296860 290310
rect 297114 290222 297294 290310
rect 297402 290222 297582 290310
rect 297690 290222 297870 290310
rect 297978 290222 298158 290310
rect 298266 290222 298446 290310
rect 298554 290222 298734 290310
rect 298842 290222 299022 290310
rect 299130 290222 299310 290310
rect 299564 290222 299744 290310
rect 299852 290222 300032 290310
rect 300140 290222 300320 290310
rect 300428 290222 300608 290310
rect 300716 290222 300896 290310
rect 301004 290222 301184 290310
rect 301292 290222 301472 290310
rect 301580 290222 301760 290310
rect 302014 290222 302194 290310
rect 302302 290222 302482 290310
rect 302590 290222 302770 290310
rect 302878 290222 303058 290310
rect 303166 290222 303346 290310
rect 303454 290222 303634 290310
rect 303742 290222 303922 290310
rect 304030 290222 304210 290310
rect 304464 290222 304644 290310
rect 304752 290222 304932 290310
rect 305040 290222 305220 290310
rect 305328 290222 305508 290310
rect 305616 290222 305796 290310
rect 305904 290222 306084 290310
rect 306192 290222 306372 290310
rect 306480 290222 306660 290310
rect 306914 290222 307094 290310
rect 307202 290222 307382 290310
rect 307490 290222 307670 290310
rect 307778 290222 307958 290310
rect 308066 290222 308246 290310
rect 308354 290222 308534 290310
rect 308642 290222 308822 290310
rect 308930 290222 309110 290310
rect 309364 290222 309544 290310
rect 309652 290222 309832 290310
rect 309940 290222 310120 290310
rect 310228 290222 310408 290310
rect 310516 290222 310696 290310
rect 310804 290222 310984 290310
rect 311092 290222 311272 290310
rect 311380 290222 311560 290310
rect 311814 290222 311994 290310
rect 312102 290222 312282 290310
rect 312390 290222 312570 290310
rect 312678 290222 312858 290310
rect 312966 290222 313146 290310
rect 313254 290222 313434 290310
rect 313542 290222 313722 290310
rect 313830 290222 314010 290310
rect 314264 290222 314444 290310
rect 314552 290222 314732 290310
rect 314840 290222 315020 290310
rect 315128 290222 315308 290310
rect 315416 290222 315596 290310
rect 315704 290222 315884 290310
rect 315992 290222 316172 290310
rect 316280 290222 316460 290310
rect 316714 290222 316894 290310
rect 317002 290222 317182 290310
rect 317290 290222 317470 290310
rect 317578 290222 317758 290310
rect 317866 290222 318046 290310
rect 318154 290222 318334 290310
rect 318442 290222 318622 290310
rect 318730 290222 318910 290310
rect 319164 290222 319344 290310
rect 319452 290222 319632 290310
rect 319740 290222 319920 290310
rect 320028 290222 320208 290310
rect 320316 290222 320496 290310
rect 320604 290222 320784 290310
rect 320892 290222 321072 290310
rect 321180 290222 321360 290310
rect 321614 290222 321794 290310
rect 321902 290222 322082 290310
rect 322190 290222 322370 290310
rect 322478 290222 322658 290310
rect 322766 290222 322946 290310
rect 323054 290222 323234 290310
rect 323342 290222 323522 290310
rect 323630 290222 323810 290310
rect 324064 290222 324244 290310
rect 324352 290222 324532 290310
rect 324640 290222 324820 290310
rect 324928 290222 325108 290310
rect 325216 290222 325396 290310
rect 325504 290222 325684 290310
rect 325792 290222 325972 290310
rect 326080 290222 326260 290310
rect 326514 290222 326694 290310
rect 326802 290222 326982 290310
rect 327090 290222 327270 290310
rect 327378 290222 327558 290310
rect 327666 290222 327846 290310
rect 327954 290222 328134 290310
rect 328242 290222 328422 290310
rect 328530 290222 328710 290310
rect 328964 290222 329144 290310
rect 329252 290222 329432 290310
rect 329540 290222 329720 290310
rect 329828 290222 330008 290310
rect 330116 290222 330296 290310
rect 330404 290222 330584 290310
rect 330692 290222 330872 290310
rect 330980 290222 331160 290310
rect 331414 290222 331594 290310
rect 331702 290222 331882 290310
rect 331990 290222 332170 290310
rect 332278 290222 332458 290310
rect 332566 290222 332746 290310
rect 332854 290222 333034 290310
rect 333142 290222 333322 290310
rect 333430 290222 333610 290310
rect 333864 290222 334044 290310
rect 334152 290222 334332 290310
rect 334440 290222 334620 290310
rect 334728 290222 334908 290310
rect 335016 290222 335196 290310
rect 335304 290222 335484 290310
rect 335592 290222 335772 290310
rect 335880 290222 336060 290310
rect 336314 290222 336494 290310
rect 336602 290222 336782 290310
rect 336890 290222 337070 290310
rect 337178 290222 337358 290310
rect 337466 290222 337646 290310
rect 337754 290222 337934 290310
rect 338042 290222 338222 290310
rect 338330 290222 338510 290310
rect 338764 290222 338944 290310
rect 339052 290222 339232 290310
rect 339340 290222 339520 290310
rect 339628 290222 339808 290310
rect 339916 290222 340096 290310
rect 340204 290222 340384 290310
rect 340492 290222 340672 290310
rect 340780 290222 340960 290310
rect 341214 290222 341394 290310
rect 341502 290222 341682 290310
rect 341790 290222 341970 290310
rect 342078 290222 342258 290310
rect 342366 290222 342546 290310
rect 342654 290222 342834 290310
rect 342942 290222 343122 290310
rect 343230 290222 343410 290310
rect 343664 290222 343844 290310
rect 343952 290222 344132 290310
rect 344240 290222 344420 290310
rect 344528 290222 344708 290310
rect 344816 290222 344996 290310
rect 345104 290222 345284 290310
rect 345392 290222 345572 290310
rect 345680 290222 345860 290310
rect 346114 290222 346294 290310
rect 346402 290222 346582 290310
rect 346690 290222 346870 290310
rect 346978 290222 347158 290310
rect 347266 290222 347446 290310
rect 347554 290222 347734 290310
rect 347842 290222 348022 290310
rect 348130 290222 348310 290310
rect 348564 290222 348744 290310
rect 348852 290222 349032 290310
rect 349140 290222 349320 290310
rect 349428 290222 349608 290310
rect 349716 290222 349896 290310
rect 350004 290222 350184 290310
rect 350292 290222 350472 290310
rect 350580 290222 350760 290310
rect 351014 290222 351194 290310
rect 351302 290222 351482 290310
rect 351590 290222 351770 290310
rect 351878 290222 352058 290310
rect 352166 290222 352346 290310
rect 352454 290222 352634 290310
rect 352742 290222 352922 290310
rect 353030 290222 353210 290310
rect 353464 290222 353644 290310
rect 353752 290222 353932 290310
rect 354040 290222 354220 290310
rect 354328 290222 354508 290310
rect 354616 290222 354796 290310
rect 354904 290222 355084 290310
rect 355192 290222 355372 290310
rect 355480 290222 355660 290310
rect 355914 290222 356094 290310
rect 356202 290222 356382 290310
rect 356490 290222 356670 290310
rect 356778 290222 356958 290310
rect 357066 290222 357246 290310
rect 357354 290222 357534 290310
rect 357642 290222 357822 290310
rect 357930 290222 358110 290310
rect 358364 290222 358544 290310
rect 358652 290222 358832 290310
rect 358940 290222 359120 290310
rect 359228 290222 359408 290310
rect 359516 290222 359696 290310
rect 359804 290222 359984 290310
rect 360092 290222 360272 290310
rect 360380 290222 360560 290310
rect 360814 290222 360994 290310
rect 361102 290222 361282 290310
rect 361390 290222 361570 290310
rect 361678 290222 361858 290310
rect 361966 290222 362146 290310
rect 362254 290222 362434 290310
rect 362542 290222 362722 290310
rect 362830 290222 363010 290310
rect 363264 290222 363444 290310
rect 363552 290222 363732 290310
rect 363840 290222 364020 290310
rect 364128 290222 364308 290310
rect 364416 290222 364596 290310
rect 364704 290222 364884 290310
rect 364992 290222 365172 290310
rect 365280 290222 365460 290310
rect 365714 290222 365894 290310
rect 366002 290222 366182 290310
rect 366290 290222 366470 290310
rect 366578 290222 366758 290310
rect 366866 290222 367046 290310
rect 367154 290222 367334 290310
rect 367442 290222 367622 290310
rect 367730 290222 367910 290310
rect 243214 290006 243394 290094
rect 243502 290006 243682 290094
rect 243790 290006 243970 290094
rect 244078 290006 244258 290094
rect 244366 290006 244546 290094
rect 244654 290006 244834 290094
rect 244942 290006 245122 290094
rect 245230 290006 245410 290094
rect 245664 290006 245844 290094
rect 245952 290006 246132 290094
rect 246240 290006 246420 290094
rect 246528 290006 246708 290094
rect 246816 290006 246996 290094
rect 247104 290006 247284 290094
rect 247392 290006 247572 290094
rect 247680 290006 247860 290094
rect 248114 290006 248294 290094
rect 248402 290006 248582 290094
rect 248690 290006 248870 290094
rect 248978 290006 249158 290094
rect 249266 290006 249446 290094
rect 249554 290006 249734 290094
rect 249842 290006 250022 290094
rect 250130 290006 250310 290094
rect 250564 290006 250744 290094
rect 250852 290006 251032 290094
rect 251140 290006 251320 290094
rect 251428 290006 251608 290094
rect 251716 290006 251896 290094
rect 252004 290006 252184 290094
rect 252292 290006 252472 290094
rect 252580 290006 252760 290094
rect 253014 290006 253194 290094
rect 253302 290006 253482 290094
rect 253590 290006 253770 290094
rect 253878 290006 254058 290094
rect 254166 290006 254346 290094
rect 254454 290006 254634 290094
rect 254742 290006 254922 290094
rect 255030 290006 255210 290094
rect 255464 290006 255644 290094
rect 255752 290006 255932 290094
rect 256040 290006 256220 290094
rect 256328 290006 256508 290094
rect 256616 290006 256796 290094
rect 256904 290006 257084 290094
rect 257192 290006 257372 290094
rect 257480 290006 257660 290094
rect 257914 290006 258094 290094
rect 258202 290006 258382 290094
rect 258490 290006 258670 290094
rect 258778 290006 258958 290094
rect 259066 290006 259246 290094
rect 259354 290006 259534 290094
rect 259642 290006 259822 290094
rect 259930 290006 260110 290094
rect 260364 290006 260544 290094
rect 260652 290006 260832 290094
rect 260940 290006 261120 290094
rect 261228 290006 261408 290094
rect 261516 290006 261696 290094
rect 261804 290006 261984 290094
rect 262092 290006 262272 290094
rect 262380 290006 262560 290094
rect 262814 290006 262994 290094
rect 263102 290006 263282 290094
rect 263390 290006 263570 290094
rect 263678 290006 263858 290094
rect 263966 290006 264146 290094
rect 264254 290006 264434 290094
rect 264542 290006 264722 290094
rect 264830 290006 265010 290094
rect 265264 290006 265444 290094
rect 265552 290006 265732 290094
rect 265840 290006 266020 290094
rect 266128 290006 266308 290094
rect 266416 290006 266596 290094
rect 266704 290006 266884 290094
rect 266992 290006 267172 290094
rect 267280 290006 267460 290094
rect 267714 290006 267894 290094
rect 268002 290006 268182 290094
rect 268290 290006 268470 290094
rect 268578 290006 268758 290094
rect 268866 290006 269046 290094
rect 269154 290006 269334 290094
rect 269442 290006 269622 290094
rect 269730 290006 269910 290094
rect 270164 290006 270344 290094
rect 270452 290006 270632 290094
rect 270740 290006 270920 290094
rect 271028 290006 271208 290094
rect 271316 290006 271496 290094
rect 271604 290006 271784 290094
rect 271892 290006 272072 290094
rect 272180 290006 272360 290094
rect 272614 290006 272794 290094
rect 272902 290006 273082 290094
rect 273190 290006 273370 290094
rect 273478 290006 273658 290094
rect 273766 290006 273946 290094
rect 274054 290006 274234 290094
rect 274342 290006 274522 290094
rect 274630 290006 274810 290094
rect 275064 290006 275244 290094
rect 275352 290006 275532 290094
rect 275640 290006 275820 290094
rect 275928 290006 276108 290094
rect 276216 290006 276396 290094
rect 276504 290006 276684 290094
rect 276792 290006 276972 290094
rect 277080 290006 277260 290094
rect 277514 290006 277694 290094
rect 277802 290006 277982 290094
rect 278090 290006 278270 290094
rect 278378 290006 278558 290094
rect 278666 290006 278846 290094
rect 278954 290006 279134 290094
rect 279242 290006 279422 290094
rect 279530 290006 279710 290094
rect 279964 290006 280144 290094
rect 280252 290006 280432 290094
rect 280540 290006 280720 290094
rect 280828 290006 281008 290094
rect 281116 290006 281296 290094
rect 281404 290006 281584 290094
rect 281692 290006 281872 290094
rect 281980 290006 282160 290094
rect 282414 290006 282594 290094
rect 282702 290006 282882 290094
rect 282990 290006 283170 290094
rect 283278 290006 283458 290094
rect 283566 290006 283746 290094
rect 283854 290006 284034 290094
rect 284142 290006 284322 290094
rect 284430 290006 284610 290094
rect 284864 290006 285044 290094
rect 285152 290006 285332 290094
rect 285440 290006 285620 290094
rect 285728 290006 285908 290094
rect 286016 290006 286196 290094
rect 286304 290006 286484 290094
rect 286592 290006 286772 290094
rect 286880 290006 287060 290094
rect 287314 290006 287494 290094
rect 287602 290006 287782 290094
rect 287890 290006 288070 290094
rect 288178 290006 288358 290094
rect 288466 290006 288646 290094
rect 288754 290006 288934 290094
rect 289042 290006 289222 290094
rect 289330 290006 289510 290094
rect 289764 290006 289944 290094
rect 290052 290006 290232 290094
rect 290340 290006 290520 290094
rect 290628 290006 290808 290094
rect 290916 290006 291096 290094
rect 291204 290006 291384 290094
rect 291492 290006 291672 290094
rect 291780 290006 291960 290094
rect 292214 290006 292394 290094
rect 292502 290006 292682 290094
rect 292790 290006 292970 290094
rect 293078 290006 293258 290094
rect 293366 290006 293546 290094
rect 293654 290006 293834 290094
rect 293942 290006 294122 290094
rect 294230 290006 294410 290094
rect 294664 290006 294844 290094
rect 294952 290006 295132 290094
rect 295240 290006 295420 290094
rect 295528 290006 295708 290094
rect 295816 290006 295996 290094
rect 296104 290006 296284 290094
rect 296392 290006 296572 290094
rect 296680 290006 296860 290094
rect 297114 290006 297294 290094
rect 297402 290006 297582 290094
rect 297690 290006 297870 290094
rect 297978 290006 298158 290094
rect 298266 290006 298446 290094
rect 298554 290006 298734 290094
rect 298842 290006 299022 290094
rect 299130 290006 299310 290094
rect 299564 290006 299744 290094
rect 299852 290006 300032 290094
rect 300140 290006 300320 290094
rect 300428 290006 300608 290094
rect 300716 290006 300896 290094
rect 301004 290006 301184 290094
rect 301292 290006 301472 290094
rect 301580 290006 301760 290094
rect 302014 290006 302194 290094
rect 302302 290006 302482 290094
rect 302590 290006 302770 290094
rect 302878 290006 303058 290094
rect 303166 290006 303346 290094
rect 303454 290006 303634 290094
rect 303742 290006 303922 290094
rect 304030 290006 304210 290094
rect 304464 290006 304644 290094
rect 304752 290006 304932 290094
rect 305040 290006 305220 290094
rect 305328 290006 305508 290094
rect 305616 290006 305796 290094
rect 305904 290006 306084 290094
rect 306192 290006 306372 290094
rect 306480 290006 306660 290094
rect 306914 290006 307094 290094
rect 307202 290006 307382 290094
rect 307490 290006 307670 290094
rect 307778 290006 307958 290094
rect 308066 290006 308246 290094
rect 308354 290006 308534 290094
rect 308642 290006 308822 290094
rect 308930 290006 309110 290094
rect 309364 290006 309544 290094
rect 309652 290006 309832 290094
rect 309940 290006 310120 290094
rect 310228 290006 310408 290094
rect 310516 290006 310696 290094
rect 310804 290006 310984 290094
rect 311092 290006 311272 290094
rect 311380 290006 311560 290094
rect 311814 290006 311994 290094
rect 312102 290006 312282 290094
rect 312390 290006 312570 290094
rect 312678 290006 312858 290094
rect 312966 290006 313146 290094
rect 313254 290006 313434 290094
rect 313542 290006 313722 290094
rect 313830 290006 314010 290094
rect 314264 290006 314444 290094
rect 314552 290006 314732 290094
rect 314840 290006 315020 290094
rect 315128 290006 315308 290094
rect 315416 290006 315596 290094
rect 315704 290006 315884 290094
rect 315992 290006 316172 290094
rect 316280 290006 316460 290094
rect 316714 290006 316894 290094
rect 317002 290006 317182 290094
rect 317290 290006 317470 290094
rect 317578 290006 317758 290094
rect 317866 290006 318046 290094
rect 318154 290006 318334 290094
rect 318442 290006 318622 290094
rect 318730 290006 318910 290094
rect 319164 290006 319344 290094
rect 319452 290006 319632 290094
rect 319740 290006 319920 290094
rect 320028 290006 320208 290094
rect 320316 290006 320496 290094
rect 320604 290006 320784 290094
rect 320892 290006 321072 290094
rect 321180 290006 321360 290094
rect 321614 290006 321794 290094
rect 321902 290006 322082 290094
rect 322190 290006 322370 290094
rect 322478 290006 322658 290094
rect 322766 290006 322946 290094
rect 323054 290006 323234 290094
rect 323342 290006 323522 290094
rect 323630 290006 323810 290094
rect 324064 290006 324244 290094
rect 324352 290006 324532 290094
rect 324640 290006 324820 290094
rect 324928 290006 325108 290094
rect 325216 290006 325396 290094
rect 325504 290006 325684 290094
rect 325792 290006 325972 290094
rect 326080 290006 326260 290094
rect 326514 290006 326694 290094
rect 326802 290006 326982 290094
rect 327090 290006 327270 290094
rect 327378 290006 327558 290094
rect 327666 290006 327846 290094
rect 327954 290006 328134 290094
rect 328242 290006 328422 290094
rect 328530 290006 328710 290094
rect 328964 290006 329144 290094
rect 329252 290006 329432 290094
rect 329540 290006 329720 290094
rect 329828 290006 330008 290094
rect 330116 290006 330296 290094
rect 330404 290006 330584 290094
rect 330692 290006 330872 290094
rect 330980 290006 331160 290094
rect 331414 290006 331594 290094
rect 331702 290006 331882 290094
rect 331990 290006 332170 290094
rect 332278 290006 332458 290094
rect 332566 290006 332746 290094
rect 332854 290006 333034 290094
rect 333142 290006 333322 290094
rect 333430 290006 333610 290094
rect 333864 290006 334044 290094
rect 334152 290006 334332 290094
rect 334440 290006 334620 290094
rect 334728 290006 334908 290094
rect 335016 290006 335196 290094
rect 335304 290006 335484 290094
rect 335592 290006 335772 290094
rect 335880 290006 336060 290094
rect 336314 290006 336494 290094
rect 336602 290006 336782 290094
rect 336890 290006 337070 290094
rect 337178 290006 337358 290094
rect 337466 290006 337646 290094
rect 337754 290006 337934 290094
rect 338042 290006 338222 290094
rect 338330 290006 338510 290094
rect 338764 290006 338944 290094
rect 339052 290006 339232 290094
rect 339340 290006 339520 290094
rect 339628 290006 339808 290094
rect 339916 290006 340096 290094
rect 340204 290006 340384 290094
rect 340492 290006 340672 290094
rect 340780 290006 340960 290094
rect 341214 290006 341394 290094
rect 341502 290006 341682 290094
rect 341790 290006 341970 290094
rect 342078 290006 342258 290094
rect 342366 290006 342546 290094
rect 342654 290006 342834 290094
rect 342942 290006 343122 290094
rect 343230 290006 343410 290094
rect 343664 290006 343844 290094
rect 343952 290006 344132 290094
rect 344240 290006 344420 290094
rect 344528 290006 344708 290094
rect 344816 290006 344996 290094
rect 345104 290006 345284 290094
rect 345392 290006 345572 290094
rect 345680 290006 345860 290094
rect 346114 290006 346294 290094
rect 346402 290006 346582 290094
rect 346690 290006 346870 290094
rect 346978 290006 347158 290094
rect 347266 290006 347446 290094
rect 347554 290006 347734 290094
rect 347842 290006 348022 290094
rect 348130 290006 348310 290094
rect 348564 290006 348744 290094
rect 348852 290006 349032 290094
rect 349140 290006 349320 290094
rect 349428 290006 349608 290094
rect 349716 290006 349896 290094
rect 350004 290006 350184 290094
rect 350292 290006 350472 290094
rect 350580 290006 350760 290094
rect 351014 290006 351194 290094
rect 351302 290006 351482 290094
rect 351590 290006 351770 290094
rect 351878 290006 352058 290094
rect 352166 290006 352346 290094
rect 352454 290006 352634 290094
rect 352742 290006 352922 290094
rect 353030 290006 353210 290094
rect 353464 290006 353644 290094
rect 353752 290006 353932 290094
rect 354040 290006 354220 290094
rect 354328 290006 354508 290094
rect 354616 290006 354796 290094
rect 354904 290006 355084 290094
rect 355192 290006 355372 290094
rect 355480 290006 355660 290094
rect 355914 290006 356094 290094
rect 356202 290006 356382 290094
rect 356490 290006 356670 290094
rect 356778 290006 356958 290094
rect 357066 290006 357246 290094
rect 357354 290006 357534 290094
rect 357642 290006 357822 290094
rect 357930 290006 358110 290094
rect 358364 290006 358544 290094
rect 358652 290006 358832 290094
rect 358940 290006 359120 290094
rect 359228 290006 359408 290094
rect 359516 290006 359696 290094
rect 359804 290006 359984 290094
rect 360092 290006 360272 290094
rect 360380 290006 360560 290094
rect 360814 290006 360994 290094
rect 361102 290006 361282 290094
rect 361390 290006 361570 290094
rect 361678 290006 361858 290094
rect 361966 290006 362146 290094
rect 362254 290006 362434 290094
rect 362542 290006 362722 290094
rect 362830 290006 363010 290094
rect 363264 290006 363444 290094
rect 363552 290006 363732 290094
rect 363840 290006 364020 290094
rect 364128 290006 364308 290094
rect 364416 290006 364596 290094
rect 364704 290006 364884 290094
rect 364992 290006 365172 290094
rect 365280 290006 365460 290094
rect 365714 290006 365894 290094
rect 366002 290006 366182 290094
rect 366290 290006 366470 290094
rect 366578 290006 366758 290094
rect 366866 290006 367046 290094
rect 367154 290006 367334 290094
rect 367442 290006 367622 290094
rect 367730 290006 367910 290094
rect 243214 289530 243394 289618
rect 243502 289530 243682 289618
rect 243790 289530 243970 289618
rect 244078 289530 244258 289618
rect 244366 289530 244546 289618
rect 244654 289530 244834 289618
rect 244942 289530 245122 289618
rect 245230 289530 245410 289618
rect 245664 289530 245844 289618
rect 245952 289530 246132 289618
rect 246240 289530 246420 289618
rect 246528 289530 246708 289618
rect 246816 289530 246996 289618
rect 247104 289530 247284 289618
rect 247392 289530 247572 289618
rect 247680 289530 247860 289618
rect 248114 289530 248294 289618
rect 248402 289530 248582 289618
rect 248690 289530 248870 289618
rect 248978 289530 249158 289618
rect 249266 289530 249446 289618
rect 249554 289530 249734 289618
rect 249842 289530 250022 289618
rect 250130 289530 250310 289618
rect 250564 289530 250744 289618
rect 250852 289530 251032 289618
rect 251140 289530 251320 289618
rect 251428 289530 251608 289618
rect 251716 289530 251896 289618
rect 252004 289530 252184 289618
rect 252292 289530 252472 289618
rect 252580 289530 252760 289618
rect 253014 289530 253194 289618
rect 253302 289530 253482 289618
rect 253590 289530 253770 289618
rect 253878 289530 254058 289618
rect 254166 289530 254346 289618
rect 254454 289530 254634 289618
rect 254742 289530 254922 289618
rect 255030 289530 255210 289618
rect 255464 289530 255644 289618
rect 255752 289530 255932 289618
rect 256040 289530 256220 289618
rect 256328 289530 256508 289618
rect 256616 289530 256796 289618
rect 256904 289530 257084 289618
rect 257192 289530 257372 289618
rect 257480 289530 257660 289618
rect 257914 289530 258094 289618
rect 258202 289530 258382 289618
rect 258490 289530 258670 289618
rect 258778 289530 258958 289618
rect 259066 289530 259246 289618
rect 259354 289530 259534 289618
rect 259642 289530 259822 289618
rect 259930 289530 260110 289618
rect 260364 289530 260544 289618
rect 260652 289530 260832 289618
rect 260940 289530 261120 289618
rect 261228 289530 261408 289618
rect 261516 289530 261696 289618
rect 261804 289530 261984 289618
rect 262092 289530 262272 289618
rect 262380 289530 262560 289618
rect 262814 289530 262994 289618
rect 263102 289530 263282 289618
rect 263390 289530 263570 289618
rect 263678 289530 263858 289618
rect 263966 289530 264146 289618
rect 264254 289530 264434 289618
rect 264542 289530 264722 289618
rect 264830 289530 265010 289618
rect 265264 289530 265444 289618
rect 265552 289530 265732 289618
rect 265840 289530 266020 289618
rect 266128 289530 266308 289618
rect 266416 289530 266596 289618
rect 266704 289530 266884 289618
rect 266992 289530 267172 289618
rect 267280 289530 267460 289618
rect 267714 289530 267894 289618
rect 268002 289530 268182 289618
rect 268290 289530 268470 289618
rect 268578 289530 268758 289618
rect 268866 289530 269046 289618
rect 269154 289530 269334 289618
rect 269442 289530 269622 289618
rect 269730 289530 269910 289618
rect 270164 289530 270344 289618
rect 270452 289530 270632 289618
rect 270740 289530 270920 289618
rect 271028 289530 271208 289618
rect 271316 289530 271496 289618
rect 271604 289530 271784 289618
rect 271892 289530 272072 289618
rect 272180 289530 272360 289618
rect 272614 289530 272794 289618
rect 272902 289530 273082 289618
rect 273190 289530 273370 289618
rect 273478 289530 273658 289618
rect 273766 289530 273946 289618
rect 274054 289530 274234 289618
rect 274342 289530 274522 289618
rect 274630 289530 274810 289618
rect 275064 289530 275244 289618
rect 275352 289530 275532 289618
rect 275640 289530 275820 289618
rect 275928 289530 276108 289618
rect 276216 289530 276396 289618
rect 276504 289530 276684 289618
rect 276792 289530 276972 289618
rect 277080 289530 277260 289618
rect 277514 289530 277694 289618
rect 277802 289530 277982 289618
rect 278090 289530 278270 289618
rect 278378 289530 278558 289618
rect 278666 289530 278846 289618
rect 278954 289530 279134 289618
rect 279242 289530 279422 289618
rect 279530 289530 279710 289618
rect 279964 289530 280144 289618
rect 280252 289530 280432 289618
rect 280540 289530 280720 289618
rect 280828 289530 281008 289618
rect 281116 289530 281296 289618
rect 281404 289530 281584 289618
rect 281692 289530 281872 289618
rect 281980 289530 282160 289618
rect 282414 289530 282594 289618
rect 282702 289530 282882 289618
rect 282990 289530 283170 289618
rect 283278 289530 283458 289618
rect 283566 289530 283746 289618
rect 283854 289530 284034 289618
rect 284142 289530 284322 289618
rect 284430 289530 284610 289618
rect 284864 289530 285044 289618
rect 285152 289530 285332 289618
rect 285440 289530 285620 289618
rect 285728 289530 285908 289618
rect 286016 289530 286196 289618
rect 286304 289530 286484 289618
rect 286592 289530 286772 289618
rect 286880 289530 287060 289618
rect 287314 289530 287494 289618
rect 287602 289530 287782 289618
rect 287890 289530 288070 289618
rect 288178 289530 288358 289618
rect 288466 289530 288646 289618
rect 288754 289530 288934 289618
rect 289042 289530 289222 289618
rect 289330 289530 289510 289618
rect 289764 289530 289944 289618
rect 290052 289530 290232 289618
rect 290340 289530 290520 289618
rect 290628 289530 290808 289618
rect 290916 289530 291096 289618
rect 291204 289530 291384 289618
rect 291492 289530 291672 289618
rect 291780 289530 291960 289618
rect 292214 289530 292394 289618
rect 292502 289530 292682 289618
rect 292790 289530 292970 289618
rect 293078 289530 293258 289618
rect 293366 289530 293546 289618
rect 293654 289530 293834 289618
rect 293942 289530 294122 289618
rect 294230 289530 294410 289618
rect 294664 289530 294844 289618
rect 294952 289530 295132 289618
rect 295240 289530 295420 289618
rect 295528 289530 295708 289618
rect 295816 289530 295996 289618
rect 296104 289530 296284 289618
rect 296392 289530 296572 289618
rect 296680 289530 296860 289618
rect 297114 289530 297294 289618
rect 297402 289530 297582 289618
rect 297690 289530 297870 289618
rect 297978 289530 298158 289618
rect 298266 289530 298446 289618
rect 298554 289530 298734 289618
rect 298842 289530 299022 289618
rect 299130 289530 299310 289618
rect 299564 289530 299744 289618
rect 299852 289530 300032 289618
rect 300140 289530 300320 289618
rect 300428 289530 300608 289618
rect 300716 289530 300896 289618
rect 301004 289530 301184 289618
rect 301292 289530 301472 289618
rect 301580 289530 301760 289618
rect 302014 289530 302194 289618
rect 302302 289530 302482 289618
rect 302590 289530 302770 289618
rect 302878 289530 303058 289618
rect 303166 289530 303346 289618
rect 303454 289530 303634 289618
rect 303742 289530 303922 289618
rect 304030 289530 304210 289618
rect 304464 289530 304644 289618
rect 304752 289530 304932 289618
rect 305040 289530 305220 289618
rect 305328 289530 305508 289618
rect 305616 289530 305796 289618
rect 305904 289530 306084 289618
rect 306192 289530 306372 289618
rect 306480 289530 306660 289618
rect 306914 289530 307094 289618
rect 307202 289530 307382 289618
rect 307490 289530 307670 289618
rect 307778 289530 307958 289618
rect 308066 289530 308246 289618
rect 308354 289530 308534 289618
rect 308642 289530 308822 289618
rect 308930 289530 309110 289618
rect 309364 289530 309544 289618
rect 309652 289530 309832 289618
rect 309940 289530 310120 289618
rect 310228 289530 310408 289618
rect 310516 289530 310696 289618
rect 310804 289530 310984 289618
rect 311092 289530 311272 289618
rect 311380 289530 311560 289618
rect 311814 289530 311994 289618
rect 312102 289530 312282 289618
rect 312390 289530 312570 289618
rect 312678 289530 312858 289618
rect 312966 289530 313146 289618
rect 313254 289530 313434 289618
rect 313542 289530 313722 289618
rect 313830 289530 314010 289618
rect 314264 289530 314444 289618
rect 314552 289530 314732 289618
rect 314840 289530 315020 289618
rect 315128 289530 315308 289618
rect 315416 289530 315596 289618
rect 315704 289530 315884 289618
rect 315992 289530 316172 289618
rect 316280 289530 316460 289618
rect 316714 289530 316894 289618
rect 317002 289530 317182 289618
rect 317290 289530 317470 289618
rect 317578 289530 317758 289618
rect 317866 289530 318046 289618
rect 318154 289530 318334 289618
rect 318442 289530 318622 289618
rect 318730 289530 318910 289618
rect 319164 289530 319344 289618
rect 319452 289530 319632 289618
rect 319740 289530 319920 289618
rect 320028 289530 320208 289618
rect 320316 289530 320496 289618
rect 320604 289530 320784 289618
rect 320892 289530 321072 289618
rect 321180 289530 321360 289618
rect 321614 289530 321794 289618
rect 321902 289530 322082 289618
rect 322190 289530 322370 289618
rect 322478 289530 322658 289618
rect 322766 289530 322946 289618
rect 323054 289530 323234 289618
rect 323342 289530 323522 289618
rect 323630 289530 323810 289618
rect 324064 289530 324244 289618
rect 324352 289530 324532 289618
rect 324640 289530 324820 289618
rect 324928 289530 325108 289618
rect 325216 289530 325396 289618
rect 325504 289530 325684 289618
rect 325792 289530 325972 289618
rect 326080 289530 326260 289618
rect 326514 289530 326694 289618
rect 326802 289530 326982 289618
rect 327090 289530 327270 289618
rect 327378 289530 327558 289618
rect 327666 289530 327846 289618
rect 327954 289530 328134 289618
rect 328242 289530 328422 289618
rect 328530 289530 328710 289618
rect 328964 289530 329144 289618
rect 329252 289530 329432 289618
rect 329540 289530 329720 289618
rect 329828 289530 330008 289618
rect 330116 289530 330296 289618
rect 330404 289530 330584 289618
rect 330692 289530 330872 289618
rect 330980 289530 331160 289618
rect 331414 289530 331594 289618
rect 331702 289530 331882 289618
rect 331990 289530 332170 289618
rect 332278 289530 332458 289618
rect 332566 289530 332746 289618
rect 332854 289530 333034 289618
rect 333142 289530 333322 289618
rect 333430 289530 333610 289618
rect 333864 289530 334044 289618
rect 334152 289530 334332 289618
rect 334440 289530 334620 289618
rect 334728 289530 334908 289618
rect 335016 289530 335196 289618
rect 335304 289530 335484 289618
rect 335592 289530 335772 289618
rect 335880 289530 336060 289618
rect 336314 289530 336494 289618
rect 336602 289530 336782 289618
rect 336890 289530 337070 289618
rect 337178 289530 337358 289618
rect 337466 289530 337646 289618
rect 337754 289530 337934 289618
rect 338042 289530 338222 289618
rect 338330 289530 338510 289618
rect 338764 289530 338944 289618
rect 339052 289530 339232 289618
rect 339340 289530 339520 289618
rect 339628 289530 339808 289618
rect 339916 289530 340096 289618
rect 340204 289530 340384 289618
rect 340492 289530 340672 289618
rect 340780 289530 340960 289618
rect 341214 289530 341394 289618
rect 341502 289530 341682 289618
rect 341790 289530 341970 289618
rect 342078 289530 342258 289618
rect 342366 289530 342546 289618
rect 342654 289530 342834 289618
rect 342942 289530 343122 289618
rect 343230 289530 343410 289618
rect 343664 289530 343844 289618
rect 343952 289530 344132 289618
rect 344240 289530 344420 289618
rect 344528 289530 344708 289618
rect 344816 289530 344996 289618
rect 345104 289530 345284 289618
rect 345392 289530 345572 289618
rect 345680 289530 345860 289618
rect 346114 289530 346294 289618
rect 346402 289530 346582 289618
rect 346690 289530 346870 289618
rect 346978 289530 347158 289618
rect 347266 289530 347446 289618
rect 347554 289530 347734 289618
rect 347842 289530 348022 289618
rect 348130 289530 348310 289618
rect 348564 289530 348744 289618
rect 348852 289530 349032 289618
rect 349140 289530 349320 289618
rect 349428 289530 349608 289618
rect 349716 289530 349896 289618
rect 350004 289530 350184 289618
rect 350292 289530 350472 289618
rect 350580 289530 350760 289618
rect 351014 289530 351194 289618
rect 351302 289530 351482 289618
rect 351590 289530 351770 289618
rect 351878 289530 352058 289618
rect 352166 289530 352346 289618
rect 352454 289530 352634 289618
rect 352742 289530 352922 289618
rect 353030 289530 353210 289618
rect 353464 289530 353644 289618
rect 353752 289530 353932 289618
rect 354040 289530 354220 289618
rect 354328 289530 354508 289618
rect 354616 289530 354796 289618
rect 354904 289530 355084 289618
rect 355192 289530 355372 289618
rect 355480 289530 355660 289618
rect 355914 289530 356094 289618
rect 356202 289530 356382 289618
rect 356490 289530 356670 289618
rect 356778 289530 356958 289618
rect 357066 289530 357246 289618
rect 357354 289530 357534 289618
rect 357642 289530 357822 289618
rect 357930 289530 358110 289618
rect 358364 289530 358544 289618
rect 358652 289530 358832 289618
rect 358940 289530 359120 289618
rect 359228 289530 359408 289618
rect 359516 289530 359696 289618
rect 359804 289530 359984 289618
rect 360092 289530 360272 289618
rect 360380 289530 360560 289618
rect 360814 289530 360994 289618
rect 361102 289530 361282 289618
rect 361390 289530 361570 289618
rect 361678 289530 361858 289618
rect 361966 289530 362146 289618
rect 362254 289530 362434 289618
rect 362542 289530 362722 289618
rect 362830 289530 363010 289618
rect 363264 289530 363444 289618
rect 363552 289530 363732 289618
rect 363840 289530 364020 289618
rect 364128 289530 364308 289618
rect 364416 289530 364596 289618
rect 364704 289530 364884 289618
rect 364992 289530 365172 289618
rect 365280 289530 365460 289618
rect 365714 289530 365894 289618
rect 366002 289530 366182 289618
rect 366290 289530 366470 289618
rect 366578 289530 366758 289618
rect 366866 289530 367046 289618
rect 367154 289530 367334 289618
rect 367442 289530 367622 289618
rect 367730 289530 367910 289618
rect 243214 289314 243394 289402
rect 243502 289314 243682 289402
rect 243790 289314 243970 289402
rect 244078 289314 244258 289402
rect 244366 289314 244546 289402
rect 244654 289314 244834 289402
rect 244942 289314 245122 289402
rect 245230 289314 245410 289402
rect 245664 289314 245844 289402
rect 245952 289314 246132 289402
rect 246240 289314 246420 289402
rect 246528 289314 246708 289402
rect 246816 289314 246996 289402
rect 247104 289314 247284 289402
rect 247392 289314 247572 289402
rect 247680 289314 247860 289402
rect 248114 289314 248294 289402
rect 248402 289314 248582 289402
rect 248690 289314 248870 289402
rect 248978 289314 249158 289402
rect 249266 289314 249446 289402
rect 249554 289314 249734 289402
rect 249842 289314 250022 289402
rect 250130 289314 250310 289402
rect 250564 289314 250744 289402
rect 360436 289314 360560 289402
rect 360814 289314 360994 289402
rect 361102 289314 361282 289402
rect 361390 289314 361570 289402
rect 361678 289314 361858 289402
rect 361966 289314 362146 289402
rect 362254 289314 362434 289402
rect 362542 289314 362722 289402
rect 362830 289314 363010 289402
rect 363264 289314 363444 289402
rect 363552 289314 363732 289402
rect 363840 289314 364020 289402
rect 364128 289314 364308 289402
rect 364416 289314 364596 289402
rect 364704 289314 364884 289402
rect 364992 289314 365172 289402
rect 365280 289314 365460 289402
rect 365714 289314 365894 289402
rect 366002 289314 366182 289402
rect 366290 289314 366470 289402
rect 366578 289314 366758 289402
rect 366866 289314 367046 289402
rect 367154 289314 367334 289402
rect 367442 289314 367622 289402
rect 367730 289314 367910 289402
rect 243214 288838 243394 288926
rect 243502 288838 243682 288926
rect 243790 288838 243970 288926
rect 244078 288838 244258 288926
rect 244366 288838 244546 288926
rect 244654 288838 244834 288926
rect 244942 288838 245122 288926
rect 245230 288838 245410 288926
rect 245664 288838 245844 288926
rect 245952 288838 246132 288926
rect 246240 288838 246420 288926
rect 246528 288838 246708 288926
rect 246816 288838 246996 288926
rect 247104 288838 247284 288926
rect 247392 288838 247572 288926
rect 247680 288838 247860 288926
rect 248114 288838 248294 288926
rect 248402 288838 248582 288926
rect 248690 288838 248870 288926
rect 248978 288838 249158 288926
rect 249266 288838 249446 288926
rect 249554 288838 249734 288926
rect 249842 288838 250022 288926
rect 250130 288838 250310 288926
rect 250564 288838 250744 288926
rect 360436 288838 360560 288926
rect 360814 288838 360994 288926
rect 361102 288838 361282 288926
rect 361390 288838 361570 288926
rect 361678 288838 361858 288926
rect 361966 288838 362146 288926
rect 362254 288838 362434 288926
rect 362542 288838 362722 288926
rect 362830 288838 363010 288926
rect 363264 288838 363444 288926
rect 363552 288838 363732 288926
rect 363840 288838 364020 288926
rect 364128 288838 364308 288926
rect 364416 288838 364596 288926
rect 364704 288838 364884 288926
rect 364992 288838 365172 288926
rect 365280 288838 365460 288926
rect 365714 288838 365894 288926
rect 366002 288838 366182 288926
rect 366290 288838 366470 288926
rect 366578 288838 366758 288926
rect 366866 288838 367046 288926
rect 367154 288838 367334 288926
rect 367442 288838 367622 288926
rect 367730 288838 367910 288926
rect 243214 288622 243394 288710
rect 243502 288622 243682 288710
rect 243790 288622 243970 288710
rect 244078 288622 244258 288710
rect 244366 288622 244546 288710
rect 244654 288622 244834 288710
rect 244942 288622 245122 288710
rect 245230 288622 245410 288710
rect 245664 288622 245844 288710
rect 245952 288622 246132 288710
rect 246240 288622 246420 288710
rect 246528 288622 246708 288710
rect 246816 288622 246996 288710
rect 247104 288622 247284 288710
rect 247392 288622 247572 288710
rect 247680 288622 247860 288710
rect 248114 288622 248294 288710
rect 248402 288622 248582 288710
rect 248690 288622 248870 288710
rect 248978 288622 249158 288710
rect 249266 288622 249446 288710
rect 249554 288622 249734 288710
rect 249842 288622 250022 288710
rect 250130 288622 250310 288710
rect 250564 288622 250744 288710
rect 360436 288622 360560 288710
rect 360814 288622 360994 288710
rect 361102 288622 361282 288710
rect 361390 288622 361570 288710
rect 361678 288622 361858 288710
rect 361966 288622 362146 288710
rect 362254 288622 362434 288710
rect 362542 288622 362722 288710
rect 362830 288622 363010 288710
rect 363264 288622 363444 288710
rect 363552 288622 363732 288710
rect 363840 288622 364020 288710
rect 364128 288622 364308 288710
rect 364416 288622 364596 288710
rect 364704 288622 364884 288710
rect 364992 288622 365172 288710
rect 365280 288622 365460 288710
rect 365714 288622 365894 288710
rect 366002 288622 366182 288710
rect 366290 288622 366470 288710
rect 366578 288622 366758 288710
rect 366866 288622 367046 288710
rect 367154 288622 367334 288710
rect 367442 288622 367622 288710
rect 367730 288622 367910 288710
rect 243214 288146 243394 288234
rect 243502 288146 243682 288234
rect 243790 288146 243970 288234
rect 244078 288146 244258 288234
rect 244366 288146 244546 288234
rect 244654 288146 244834 288234
rect 244942 288146 245122 288234
rect 245230 288146 245410 288234
rect 245664 288146 245844 288234
rect 245952 288146 246132 288234
rect 246240 288146 246420 288234
rect 246528 288146 246708 288234
rect 246816 288146 246996 288234
rect 247104 288146 247284 288234
rect 247392 288146 247572 288234
rect 247680 288146 247860 288234
rect 248114 288146 248294 288234
rect 248402 288146 248582 288234
rect 248690 288146 248870 288234
rect 248978 288146 249158 288234
rect 249266 288146 249446 288234
rect 249554 288146 249734 288234
rect 249842 288146 250022 288234
rect 250130 288146 250310 288234
rect 250564 288146 250744 288234
rect 360436 288146 360560 288234
rect 360814 288146 360994 288234
rect 361102 288146 361282 288234
rect 361390 288146 361570 288234
rect 361678 288146 361858 288234
rect 361966 288146 362146 288234
rect 362254 288146 362434 288234
rect 362542 288146 362722 288234
rect 362830 288146 363010 288234
rect 363264 288146 363444 288234
rect 363552 288146 363732 288234
rect 363840 288146 364020 288234
rect 364128 288146 364308 288234
rect 364416 288146 364596 288234
rect 364704 288146 364884 288234
rect 364992 288146 365172 288234
rect 365280 288146 365460 288234
rect 365714 288146 365894 288234
rect 366002 288146 366182 288234
rect 366290 288146 366470 288234
rect 366578 288146 366758 288234
rect 366866 288146 367046 288234
rect 367154 288146 367334 288234
rect 367442 288146 367622 288234
rect 367730 288146 367910 288234
rect 243214 287672 243394 287760
rect 243502 287672 243682 287760
rect 243790 287672 243970 287760
rect 244078 287672 244258 287760
rect 244366 287672 244546 287760
rect 244654 287672 244834 287760
rect 244942 287672 245122 287760
rect 245230 287672 245410 287760
rect 245664 287672 245844 287760
rect 245952 287672 246132 287760
rect 246240 287672 246420 287760
rect 246528 287672 246708 287760
rect 246816 287672 246996 287760
rect 247104 287672 247284 287760
rect 247392 287672 247572 287760
rect 247680 287672 247860 287760
rect 248114 287672 248294 287760
rect 248402 287672 248582 287760
rect 248690 287672 248870 287760
rect 248978 287672 249158 287760
rect 249266 287672 249446 287760
rect 249554 287672 249734 287760
rect 249842 287672 250022 287760
rect 250130 287672 250310 287760
rect 250564 287672 250744 287760
rect 360436 287672 360560 287760
rect 360814 287672 360994 287760
rect 361102 287672 361282 287760
rect 361390 287672 361570 287760
rect 361678 287672 361858 287760
rect 361966 287672 362146 287760
rect 362254 287672 362434 287760
rect 362542 287672 362722 287760
rect 362830 287672 363010 287760
rect 363264 287672 363444 287760
rect 363552 287672 363732 287760
rect 363840 287672 364020 287760
rect 364128 287672 364308 287760
rect 364416 287672 364596 287760
rect 364704 287672 364884 287760
rect 364992 287672 365172 287760
rect 365280 287672 365460 287760
rect 365714 287672 365894 287760
rect 366002 287672 366182 287760
rect 366290 287672 366470 287760
rect 366578 287672 366758 287760
rect 366866 287672 367046 287760
rect 367154 287672 367334 287760
rect 367442 287672 367622 287760
rect 367730 287672 367910 287760
rect 243214 287196 243394 287284
rect 243502 287196 243682 287284
rect 243790 287196 243970 287284
rect 244078 287196 244258 287284
rect 244366 287196 244546 287284
rect 244654 287196 244834 287284
rect 244942 287196 245122 287284
rect 245230 287196 245410 287284
rect 245664 287196 245844 287284
rect 245952 287196 246132 287284
rect 246240 287196 246420 287284
rect 246528 287196 246708 287284
rect 246816 287196 246996 287284
rect 247104 287196 247284 287284
rect 247392 287196 247572 287284
rect 247680 287196 247860 287284
rect 248114 287196 248294 287284
rect 248402 287196 248582 287284
rect 248690 287196 248870 287284
rect 248978 287196 249158 287284
rect 249266 287196 249446 287284
rect 249554 287196 249734 287284
rect 249842 287196 250022 287284
rect 250130 287196 250310 287284
rect 250564 287196 250744 287284
rect 360436 287196 360560 287284
rect 360814 287196 360994 287284
rect 361102 287196 361282 287284
rect 361390 287196 361570 287284
rect 361678 287196 361858 287284
rect 361966 287196 362146 287284
rect 362254 287196 362434 287284
rect 362542 287196 362722 287284
rect 362830 287196 363010 287284
rect 363264 287196 363444 287284
rect 363552 287196 363732 287284
rect 363840 287196 364020 287284
rect 364128 287196 364308 287284
rect 364416 287196 364596 287284
rect 364704 287196 364884 287284
rect 364992 287196 365172 287284
rect 365280 287196 365460 287284
rect 365714 287196 365894 287284
rect 366002 287196 366182 287284
rect 366290 287196 366470 287284
rect 366578 287196 366758 287284
rect 366866 287196 367046 287284
rect 367154 287196 367334 287284
rect 367442 287196 367622 287284
rect 367730 287196 367910 287284
rect 243214 286980 243394 287068
rect 243502 286980 243682 287068
rect 243790 286980 243970 287068
rect 244078 286980 244258 287068
rect 244366 286980 244546 287068
rect 244654 286980 244834 287068
rect 244942 286980 245122 287068
rect 245230 286980 245410 287068
rect 245664 286980 245844 287068
rect 245952 286980 246132 287068
rect 246240 286980 246420 287068
rect 246528 286980 246708 287068
rect 246816 286980 246996 287068
rect 247104 286980 247284 287068
rect 247392 286980 247572 287068
rect 247680 286980 247860 287068
rect 248114 286980 248294 287068
rect 248402 286980 248582 287068
rect 248690 286980 248870 287068
rect 248978 286980 249158 287068
rect 249266 286980 249446 287068
rect 249554 286980 249734 287068
rect 249842 286980 250022 287068
rect 250130 286980 250310 287068
rect 250564 286980 250744 287068
rect 360436 286980 360560 287068
rect 360814 286980 360994 287068
rect 361102 286980 361282 287068
rect 361390 286980 361570 287068
rect 361678 286980 361858 287068
rect 361966 286980 362146 287068
rect 362254 286980 362434 287068
rect 362542 286980 362722 287068
rect 362830 286980 363010 287068
rect 363264 286980 363444 287068
rect 363552 286980 363732 287068
rect 363840 286980 364020 287068
rect 364128 286980 364308 287068
rect 364416 286980 364596 287068
rect 364704 286980 364884 287068
rect 364992 286980 365172 287068
rect 365280 286980 365460 287068
rect 365714 286980 365894 287068
rect 366002 286980 366182 287068
rect 366290 286980 366470 287068
rect 366578 286980 366758 287068
rect 366866 286980 367046 287068
rect 367154 286980 367334 287068
rect 367442 286980 367622 287068
rect 367730 286980 367910 287068
rect 243214 286504 243394 286592
rect 243502 286504 243682 286592
rect 243790 286504 243970 286592
rect 244078 286504 244258 286592
rect 244366 286504 244546 286592
rect 244654 286504 244834 286592
rect 244942 286504 245122 286592
rect 245230 286504 245410 286592
rect 245664 286504 245844 286592
rect 245952 286504 246132 286592
rect 246240 286504 246420 286592
rect 246528 286504 246708 286592
rect 246816 286504 246996 286592
rect 247104 286504 247284 286592
rect 247392 286504 247572 286592
rect 247680 286504 247860 286592
rect 248114 286504 248294 286592
rect 248402 286504 248582 286592
rect 248690 286504 248870 286592
rect 248978 286504 249158 286592
rect 249266 286504 249446 286592
rect 249554 286504 249734 286592
rect 249842 286504 250022 286592
rect 250130 286504 250310 286592
rect 250564 286504 250744 286592
rect 360436 286504 360560 286592
rect 360814 286504 360994 286592
rect 361102 286504 361282 286592
rect 361390 286504 361570 286592
rect 361678 286504 361858 286592
rect 361966 286504 362146 286592
rect 362254 286504 362434 286592
rect 362542 286504 362722 286592
rect 362830 286504 363010 286592
rect 363264 286504 363444 286592
rect 363552 286504 363732 286592
rect 363840 286504 364020 286592
rect 364128 286504 364308 286592
rect 364416 286504 364596 286592
rect 364704 286504 364884 286592
rect 364992 286504 365172 286592
rect 365280 286504 365460 286592
rect 365714 286504 365894 286592
rect 366002 286504 366182 286592
rect 366290 286504 366470 286592
rect 366578 286504 366758 286592
rect 366866 286504 367046 286592
rect 367154 286504 367334 286592
rect 367442 286504 367622 286592
rect 367730 286504 367910 286592
rect 243214 286288 243394 286376
rect 243502 286288 243682 286376
rect 243790 286288 243970 286376
rect 244078 286288 244258 286376
rect 244366 286288 244546 286376
rect 244654 286288 244834 286376
rect 244942 286288 245122 286376
rect 245230 286288 245410 286376
rect 245664 286288 245844 286376
rect 245952 286288 246132 286376
rect 246240 286288 246420 286376
rect 246528 286288 246708 286376
rect 246816 286288 246996 286376
rect 247104 286288 247284 286376
rect 247392 286288 247572 286376
rect 247680 286288 247860 286376
rect 248114 286288 248294 286376
rect 248402 286288 248582 286376
rect 248690 286288 248870 286376
rect 248978 286288 249158 286376
rect 249266 286288 249446 286376
rect 249554 286288 249734 286376
rect 249842 286288 250022 286376
rect 250130 286288 250310 286376
rect 250564 286288 250744 286376
rect 360436 286288 360560 286376
rect 360814 286288 360994 286376
rect 361102 286288 361282 286376
rect 361390 286288 361570 286376
rect 361678 286288 361858 286376
rect 361966 286288 362146 286376
rect 362254 286288 362434 286376
rect 362542 286288 362722 286376
rect 362830 286288 363010 286376
rect 363264 286288 363444 286376
rect 363552 286288 363732 286376
rect 363840 286288 364020 286376
rect 364128 286288 364308 286376
rect 364416 286288 364596 286376
rect 364704 286288 364884 286376
rect 364992 286288 365172 286376
rect 365280 286288 365460 286376
rect 365714 286288 365894 286376
rect 366002 286288 366182 286376
rect 366290 286288 366470 286376
rect 366578 286288 366758 286376
rect 366866 286288 367046 286376
rect 367154 286288 367334 286376
rect 367442 286288 367622 286376
rect 367730 286288 367910 286376
rect 243214 285812 243394 285900
rect 243502 285812 243682 285900
rect 243790 285812 243970 285900
rect 244078 285812 244258 285900
rect 244366 285812 244546 285900
rect 244654 285812 244834 285900
rect 244942 285812 245122 285900
rect 245230 285812 245410 285900
rect 245664 285812 245844 285900
rect 245952 285812 246132 285900
rect 246240 285812 246420 285900
rect 246528 285812 246708 285900
rect 246816 285812 246996 285900
rect 247104 285812 247284 285900
rect 247392 285812 247572 285900
rect 247680 285812 247860 285900
rect 248114 285812 248294 285900
rect 248402 285812 248582 285900
rect 248690 285812 248870 285900
rect 248978 285812 249158 285900
rect 249266 285812 249446 285900
rect 249554 285812 249734 285900
rect 249842 285812 250022 285900
rect 250130 285812 250310 285900
rect 250564 285812 250744 285900
rect 360436 285812 360560 285900
rect 360814 285812 360994 285900
rect 361102 285812 361282 285900
rect 361390 285812 361570 285900
rect 361678 285812 361858 285900
rect 361966 285812 362146 285900
rect 362254 285812 362434 285900
rect 362542 285812 362722 285900
rect 362830 285812 363010 285900
rect 363264 285812 363444 285900
rect 363552 285812 363732 285900
rect 363840 285812 364020 285900
rect 364128 285812 364308 285900
rect 364416 285812 364596 285900
rect 364704 285812 364884 285900
rect 364992 285812 365172 285900
rect 365280 285812 365460 285900
rect 365714 285812 365894 285900
rect 366002 285812 366182 285900
rect 366290 285812 366470 285900
rect 366578 285812 366758 285900
rect 366866 285812 367046 285900
rect 367154 285812 367334 285900
rect 367442 285812 367622 285900
rect 367730 285812 367910 285900
rect 243214 285596 243394 285684
rect 243502 285596 243682 285684
rect 243790 285596 243970 285684
rect 244078 285596 244258 285684
rect 244366 285596 244546 285684
rect 244654 285596 244834 285684
rect 244942 285596 245122 285684
rect 245230 285596 245410 285684
rect 245664 285596 245844 285684
rect 245952 285596 246132 285684
rect 246240 285596 246420 285684
rect 246528 285596 246708 285684
rect 246816 285596 246996 285684
rect 247104 285596 247284 285684
rect 247392 285596 247572 285684
rect 247680 285596 247860 285684
rect 248114 285596 248294 285684
rect 248402 285596 248582 285684
rect 248690 285596 248870 285684
rect 248978 285596 249158 285684
rect 249266 285596 249446 285684
rect 249554 285596 249734 285684
rect 249842 285596 250022 285684
rect 250130 285596 250310 285684
rect 250564 285596 250744 285684
rect 360436 285596 360560 285684
rect 360814 285596 360994 285684
rect 361102 285596 361282 285684
rect 361390 285596 361570 285684
rect 361678 285596 361858 285684
rect 361966 285596 362146 285684
rect 362254 285596 362434 285684
rect 362542 285596 362722 285684
rect 362830 285596 363010 285684
rect 363264 285596 363444 285684
rect 363552 285596 363732 285684
rect 363840 285596 364020 285684
rect 364128 285596 364308 285684
rect 364416 285596 364596 285684
rect 364704 285596 364884 285684
rect 364992 285596 365172 285684
rect 365280 285596 365460 285684
rect 365714 285596 365894 285684
rect 366002 285596 366182 285684
rect 366290 285596 366470 285684
rect 366578 285596 366758 285684
rect 366866 285596 367046 285684
rect 367154 285596 367334 285684
rect 367442 285596 367622 285684
rect 367730 285596 367910 285684
rect 243214 285120 243394 285208
rect 243502 285120 243682 285208
rect 243790 285120 243970 285208
rect 244078 285120 244258 285208
rect 244366 285120 244546 285208
rect 244654 285120 244834 285208
rect 244942 285120 245122 285208
rect 245230 285120 245410 285208
rect 245664 285120 245844 285208
rect 245952 285120 246132 285208
rect 246240 285120 246420 285208
rect 246528 285120 246708 285208
rect 246816 285120 246996 285208
rect 247104 285120 247284 285208
rect 247392 285120 247572 285208
rect 247680 285120 247860 285208
rect 248114 285120 248294 285208
rect 248402 285120 248582 285208
rect 248690 285120 248870 285208
rect 248978 285120 249158 285208
rect 249266 285120 249446 285208
rect 249554 285120 249734 285208
rect 249842 285120 250022 285208
rect 250130 285120 250310 285208
rect 250564 285120 250744 285208
rect 360436 285120 360560 285208
rect 360814 285120 360994 285208
rect 361102 285120 361282 285208
rect 361390 285120 361570 285208
rect 361678 285120 361858 285208
rect 361966 285120 362146 285208
rect 362254 285120 362434 285208
rect 362542 285120 362722 285208
rect 362830 285120 363010 285208
rect 363264 285120 363444 285208
rect 363552 285120 363732 285208
rect 363840 285120 364020 285208
rect 364128 285120 364308 285208
rect 364416 285120 364596 285208
rect 364704 285120 364884 285208
rect 364992 285120 365172 285208
rect 365280 285120 365460 285208
rect 365714 285120 365894 285208
rect 366002 285120 366182 285208
rect 366290 285120 366470 285208
rect 366578 285120 366758 285208
rect 366866 285120 367046 285208
rect 367154 285120 367334 285208
rect 367442 285120 367622 285208
rect 367730 285120 367910 285208
rect 243214 284646 243394 284734
rect 243502 284646 243682 284734
rect 243790 284646 243970 284734
rect 244078 284646 244258 284734
rect 244366 284646 244546 284734
rect 244654 284646 244834 284734
rect 244942 284646 245122 284734
rect 245230 284646 245410 284734
rect 245664 284646 245844 284734
rect 245952 284646 246132 284734
rect 246240 284646 246420 284734
rect 246528 284646 246708 284734
rect 246816 284646 246996 284734
rect 247104 284646 247284 284734
rect 247392 284646 247572 284734
rect 247680 284646 247860 284734
rect 248114 284646 248294 284734
rect 248402 284646 248582 284734
rect 248690 284646 248870 284734
rect 248978 284646 249158 284734
rect 249266 284646 249446 284734
rect 249554 284646 249734 284734
rect 249842 284646 250022 284734
rect 250130 284646 250310 284734
rect 250564 284646 250744 284734
rect 360436 284646 360560 284734
rect 360814 284646 360994 284734
rect 361102 284646 361282 284734
rect 361390 284646 361570 284734
rect 361678 284646 361858 284734
rect 361966 284646 362146 284734
rect 362254 284646 362434 284734
rect 362542 284646 362722 284734
rect 362830 284646 363010 284734
rect 363264 284646 363444 284734
rect 363552 284646 363732 284734
rect 363840 284646 364020 284734
rect 364128 284646 364308 284734
rect 364416 284646 364596 284734
rect 364704 284646 364884 284734
rect 364992 284646 365172 284734
rect 365280 284646 365460 284734
rect 365714 284646 365894 284734
rect 366002 284646 366182 284734
rect 366290 284646 366470 284734
rect 366578 284646 366758 284734
rect 366866 284646 367046 284734
rect 367154 284646 367334 284734
rect 367442 284646 367622 284734
rect 367730 284646 367910 284734
rect 243214 284170 243394 284258
rect 243502 284170 243682 284258
rect 243790 284170 243970 284258
rect 244078 284170 244258 284258
rect 244366 284170 244546 284258
rect 244654 284170 244834 284258
rect 244942 284170 245122 284258
rect 245230 284170 245410 284258
rect 245664 284170 245844 284258
rect 245952 284170 246132 284258
rect 246240 284170 246420 284258
rect 246528 284170 246708 284258
rect 246816 284170 246996 284258
rect 247104 284170 247284 284258
rect 247392 284170 247572 284258
rect 247680 284170 247860 284258
rect 248114 284170 248294 284258
rect 248402 284170 248582 284258
rect 248690 284170 248870 284258
rect 248978 284170 249158 284258
rect 249266 284170 249446 284258
rect 249554 284170 249734 284258
rect 249842 284170 250022 284258
rect 250130 284170 250310 284258
rect 250564 284170 250744 284258
rect 360436 284170 360560 284258
rect 360814 284170 360994 284258
rect 361102 284170 361282 284258
rect 361390 284170 361570 284258
rect 361678 284170 361858 284258
rect 361966 284170 362146 284258
rect 362254 284170 362434 284258
rect 362542 284170 362722 284258
rect 362830 284170 363010 284258
rect 363264 284170 363444 284258
rect 363552 284170 363732 284258
rect 363840 284170 364020 284258
rect 364128 284170 364308 284258
rect 364416 284170 364596 284258
rect 364704 284170 364884 284258
rect 364992 284170 365172 284258
rect 365280 284170 365460 284258
rect 365714 284170 365894 284258
rect 366002 284170 366182 284258
rect 366290 284170 366470 284258
rect 366578 284170 366758 284258
rect 366866 284170 367046 284258
rect 367154 284170 367334 284258
rect 367442 284170 367622 284258
rect 367730 284170 367910 284258
rect 243214 283954 243394 284042
rect 243502 283954 243682 284042
rect 243790 283954 243970 284042
rect 244078 283954 244258 284042
rect 244366 283954 244546 284042
rect 244654 283954 244834 284042
rect 244942 283954 245122 284042
rect 245230 283954 245410 284042
rect 245664 283954 245844 284042
rect 245952 283954 246132 284042
rect 246240 283954 246420 284042
rect 246528 283954 246708 284042
rect 246816 283954 246996 284042
rect 247104 283954 247284 284042
rect 247392 283954 247572 284042
rect 247680 283954 247860 284042
rect 248114 283954 248294 284042
rect 248402 283954 248582 284042
rect 248690 283954 248870 284042
rect 248978 283954 249158 284042
rect 249266 283954 249446 284042
rect 249554 283954 249734 284042
rect 249842 283954 250022 284042
rect 250130 283954 250310 284042
rect 250564 283954 250744 284042
rect 360436 283954 360560 284042
rect 360814 283954 360994 284042
rect 361102 283954 361282 284042
rect 361390 283954 361570 284042
rect 361678 283954 361858 284042
rect 361966 283954 362146 284042
rect 362254 283954 362434 284042
rect 362542 283954 362722 284042
rect 362830 283954 363010 284042
rect 363264 283954 363444 284042
rect 363552 283954 363732 284042
rect 363840 283954 364020 284042
rect 364128 283954 364308 284042
rect 364416 283954 364596 284042
rect 364704 283954 364884 284042
rect 364992 283954 365172 284042
rect 365280 283954 365460 284042
rect 365714 283954 365894 284042
rect 366002 283954 366182 284042
rect 366290 283954 366470 284042
rect 366578 283954 366758 284042
rect 366866 283954 367046 284042
rect 367154 283954 367334 284042
rect 367442 283954 367622 284042
rect 367730 283954 367910 284042
rect 243214 283478 243394 283566
rect 243502 283478 243682 283566
rect 243790 283478 243970 283566
rect 244078 283478 244258 283566
rect 244366 283478 244546 283566
rect 244654 283478 244834 283566
rect 244942 283478 245122 283566
rect 245230 283478 245410 283566
rect 245664 283478 245844 283566
rect 245952 283478 246132 283566
rect 246240 283478 246420 283566
rect 246528 283478 246708 283566
rect 246816 283478 246996 283566
rect 247104 283478 247284 283566
rect 247392 283478 247572 283566
rect 247680 283478 247860 283566
rect 248114 283478 248294 283566
rect 248402 283478 248582 283566
rect 248690 283478 248870 283566
rect 248978 283478 249158 283566
rect 249266 283478 249446 283566
rect 249554 283478 249734 283566
rect 249842 283478 250022 283566
rect 250130 283478 250310 283566
rect 250564 283478 250744 283566
rect 360436 283478 360560 283566
rect 360814 283478 360994 283566
rect 361102 283478 361282 283566
rect 361390 283478 361570 283566
rect 361678 283478 361858 283566
rect 361966 283478 362146 283566
rect 362254 283478 362434 283566
rect 362542 283478 362722 283566
rect 362830 283478 363010 283566
rect 363264 283478 363444 283566
rect 363552 283478 363732 283566
rect 363840 283478 364020 283566
rect 364128 283478 364308 283566
rect 364416 283478 364596 283566
rect 364704 283478 364884 283566
rect 364992 283478 365172 283566
rect 365280 283478 365460 283566
rect 365714 283478 365894 283566
rect 366002 283478 366182 283566
rect 366290 283478 366470 283566
rect 366578 283478 366758 283566
rect 366866 283478 367046 283566
rect 367154 283478 367334 283566
rect 367442 283478 367622 283566
rect 367730 283478 367910 283566
rect 243214 283262 243394 283350
rect 243502 283262 243682 283350
rect 243790 283262 243970 283350
rect 244078 283262 244258 283350
rect 244366 283262 244546 283350
rect 244654 283262 244834 283350
rect 244942 283262 245122 283350
rect 245230 283262 245410 283350
rect 245664 283262 245844 283350
rect 245952 283262 246132 283350
rect 246240 283262 246420 283350
rect 246528 283262 246708 283350
rect 246816 283262 246996 283350
rect 247104 283262 247284 283350
rect 247392 283262 247572 283350
rect 247680 283262 247860 283350
rect 248114 283262 248294 283350
rect 248402 283262 248582 283350
rect 248690 283262 248870 283350
rect 248978 283262 249158 283350
rect 249266 283262 249446 283350
rect 249554 283262 249734 283350
rect 249842 283262 250022 283350
rect 250130 283262 250310 283350
rect 250564 283262 250744 283350
rect 360436 283262 360560 283350
rect 360814 283262 360994 283350
rect 361102 283262 361282 283350
rect 361390 283262 361570 283350
rect 361678 283262 361858 283350
rect 361966 283262 362146 283350
rect 362254 283262 362434 283350
rect 362542 283262 362722 283350
rect 362830 283262 363010 283350
rect 363264 283262 363444 283350
rect 363552 283262 363732 283350
rect 363840 283262 364020 283350
rect 364128 283262 364308 283350
rect 364416 283262 364596 283350
rect 364704 283262 364884 283350
rect 364992 283262 365172 283350
rect 365280 283262 365460 283350
rect 365714 283262 365894 283350
rect 366002 283262 366182 283350
rect 366290 283262 366470 283350
rect 366578 283262 366758 283350
rect 366866 283262 367046 283350
rect 367154 283262 367334 283350
rect 367442 283262 367622 283350
rect 367730 283262 367910 283350
rect 243214 282786 243394 282874
rect 243502 282786 243682 282874
rect 243790 282786 243970 282874
rect 244078 282786 244258 282874
rect 244366 282786 244546 282874
rect 244654 282786 244834 282874
rect 244942 282786 245122 282874
rect 245230 282786 245410 282874
rect 245664 282786 245844 282874
rect 245952 282786 246132 282874
rect 246240 282786 246420 282874
rect 246528 282786 246708 282874
rect 246816 282786 246996 282874
rect 247104 282786 247284 282874
rect 247392 282786 247572 282874
rect 247680 282786 247860 282874
rect 248114 282786 248294 282874
rect 248402 282786 248582 282874
rect 248690 282786 248870 282874
rect 248978 282786 249158 282874
rect 249266 282786 249446 282874
rect 249554 282786 249734 282874
rect 249842 282786 250022 282874
rect 250130 282786 250310 282874
rect 250564 282786 250744 282874
rect 360436 282786 360560 282874
rect 360814 282786 360994 282874
rect 361102 282786 361282 282874
rect 361390 282786 361570 282874
rect 361678 282786 361858 282874
rect 361966 282786 362146 282874
rect 362254 282786 362434 282874
rect 362542 282786 362722 282874
rect 362830 282786 363010 282874
rect 363264 282786 363444 282874
rect 363552 282786 363732 282874
rect 363840 282786 364020 282874
rect 364128 282786 364308 282874
rect 364416 282786 364596 282874
rect 364704 282786 364884 282874
rect 364992 282786 365172 282874
rect 365280 282786 365460 282874
rect 365714 282786 365894 282874
rect 366002 282786 366182 282874
rect 366290 282786 366470 282874
rect 366578 282786 366758 282874
rect 366866 282786 367046 282874
rect 367154 282786 367334 282874
rect 367442 282786 367622 282874
rect 367730 282786 367910 282874
rect 243214 282570 243394 282658
rect 243502 282570 243682 282658
rect 243790 282570 243970 282658
rect 244078 282570 244258 282658
rect 244366 282570 244546 282658
rect 244654 282570 244834 282658
rect 244942 282570 245122 282658
rect 245230 282570 245410 282658
rect 245664 282570 245844 282658
rect 245952 282570 246132 282658
rect 246240 282570 246420 282658
rect 246528 282570 246708 282658
rect 246816 282570 246996 282658
rect 247104 282570 247284 282658
rect 247392 282570 247572 282658
rect 247680 282570 247860 282658
rect 248114 282570 248294 282658
rect 248402 282570 248582 282658
rect 248690 282570 248870 282658
rect 248978 282570 249158 282658
rect 249266 282570 249446 282658
rect 249554 282570 249734 282658
rect 249842 282570 250022 282658
rect 250130 282570 250310 282658
rect 250564 282570 250744 282658
rect 360436 282570 360560 282658
rect 360814 282570 360994 282658
rect 361102 282570 361282 282658
rect 361390 282570 361570 282658
rect 361678 282570 361858 282658
rect 361966 282570 362146 282658
rect 362254 282570 362434 282658
rect 362542 282570 362722 282658
rect 362830 282570 363010 282658
rect 363264 282570 363444 282658
rect 363552 282570 363732 282658
rect 363840 282570 364020 282658
rect 364128 282570 364308 282658
rect 364416 282570 364596 282658
rect 364704 282570 364884 282658
rect 364992 282570 365172 282658
rect 365280 282570 365460 282658
rect 365714 282570 365894 282658
rect 366002 282570 366182 282658
rect 366290 282570 366470 282658
rect 366578 282570 366758 282658
rect 366866 282570 367046 282658
rect 367154 282570 367334 282658
rect 367442 282570 367622 282658
rect 367730 282570 367910 282658
rect 243214 282094 243394 282182
rect 243502 282094 243682 282182
rect 243790 282094 243970 282182
rect 244078 282094 244258 282182
rect 244366 282094 244546 282182
rect 244654 282094 244834 282182
rect 244942 282094 245122 282182
rect 245230 282094 245410 282182
rect 245664 282094 245844 282182
rect 245952 282094 246132 282182
rect 246240 282094 246420 282182
rect 246528 282094 246708 282182
rect 246816 282094 246996 282182
rect 247104 282094 247284 282182
rect 247392 282094 247572 282182
rect 247680 282094 247860 282182
rect 248114 282094 248294 282182
rect 248402 282094 248582 282182
rect 248690 282094 248870 282182
rect 248978 282094 249158 282182
rect 249266 282094 249446 282182
rect 249554 282094 249734 282182
rect 249842 282094 250022 282182
rect 250130 282094 250310 282182
rect 250564 282094 250744 282182
rect 360436 282094 360560 282182
rect 360814 282094 360994 282182
rect 361102 282094 361282 282182
rect 361390 282094 361570 282182
rect 361678 282094 361858 282182
rect 361966 282094 362146 282182
rect 362254 282094 362434 282182
rect 362542 282094 362722 282182
rect 362830 282094 363010 282182
rect 363264 282094 363444 282182
rect 363552 282094 363732 282182
rect 363840 282094 364020 282182
rect 364128 282094 364308 282182
rect 364416 282094 364596 282182
rect 364704 282094 364884 282182
rect 364992 282094 365172 282182
rect 365280 282094 365460 282182
rect 365714 282094 365894 282182
rect 366002 282094 366182 282182
rect 366290 282094 366470 282182
rect 366578 282094 366758 282182
rect 366866 282094 367046 282182
rect 367154 282094 367334 282182
rect 367442 282094 367622 282182
rect 367730 282094 367910 282182
rect 243214 281620 243394 281708
rect 243502 281620 243682 281708
rect 243790 281620 243970 281708
rect 244078 281620 244258 281708
rect 244366 281620 244546 281708
rect 244654 281620 244834 281708
rect 244942 281620 245122 281708
rect 245230 281620 245410 281708
rect 245664 281620 245844 281708
rect 245952 281620 246132 281708
rect 246240 281620 246420 281708
rect 246528 281620 246708 281708
rect 246816 281620 246996 281708
rect 247104 281620 247284 281708
rect 247392 281620 247572 281708
rect 247680 281620 247860 281708
rect 248114 281620 248294 281708
rect 248402 281620 248582 281708
rect 248690 281620 248870 281708
rect 248978 281620 249158 281708
rect 249266 281620 249446 281708
rect 249554 281620 249734 281708
rect 249842 281620 250022 281708
rect 250130 281620 250310 281708
rect 250564 281620 250744 281708
rect 360436 281620 360560 281708
rect 360814 281620 360994 281708
rect 361102 281620 361282 281708
rect 361390 281620 361570 281708
rect 361678 281620 361858 281708
rect 361966 281620 362146 281708
rect 362254 281620 362434 281708
rect 362542 281620 362722 281708
rect 362830 281620 363010 281708
rect 363264 281620 363444 281708
rect 363552 281620 363732 281708
rect 363840 281620 364020 281708
rect 364128 281620 364308 281708
rect 364416 281620 364596 281708
rect 364704 281620 364884 281708
rect 364992 281620 365172 281708
rect 365280 281620 365460 281708
rect 365714 281620 365894 281708
rect 366002 281620 366182 281708
rect 366290 281620 366470 281708
rect 366578 281620 366758 281708
rect 366866 281620 367046 281708
rect 367154 281620 367334 281708
rect 367442 281620 367622 281708
rect 367730 281620 367910 281708
rect 243214 281144 243394 281232
rect 243502 281144 243682 281232
rect 243790 281144 243970 281232
rect 244078 281144 244258 281232
rect 244366 281144 244546 281232
rect 244654 281144 244834 281232
rect 244942 281144 245122 281232
rect 245230 281144 245410 281232
rect 245664 281144 245844 281232
rect 245952 281144 246132 281232
rect 246240 281144 246420 281232
rect 246528 281144 246708 281232
rect 246816 281144 246996 281232
rect 247104 281144 247284 281232
rect 247392 281144 247572 281232
rect 247680 281144 247860 281232
rect 248114 281144 248294 281232
rect 248402 281144 248582 281232
rect 248690 281144 248870 281232
rect 248978 281144 249158 281232
rect 249266 281144 249446 281232
rect 249554 281144 249734 281232
rect 249842 281144 250022 281232
rect 250130 281144 250310 281232
rect 250564 281144 250744 281232
rect 360436 281144 360560 281232
rect 360814 281144 360994 281232
rect 361102 281144 361282 281232
rect 361390 281144 361570 281232
rect 361678 281144 361858 281232
rect 361966 281144 362146 281232
rect 362254 281144 362434 281232
rect 362542 281144 362722 281232
rect 362830 281144 363010 281232
rect 363264 281144 363444 281232
rect 363552 281144 363732 281232
rect 363840 281144 364020 281232
rect 364128 281144 364308 281232
rect 364416 281144 364596 281232
rect 364704 281144 364884 281232
rect 364992 281144 365172 281232
rect 365280 281144 365460 281232
rect 365714 281144 365894 281232
rect 366002 281144 366182 281232
rect 366290 281144 366470 281232
rect 366578 281144 366758 281232
rect 366866 281144 367046 281232
rect 367154 281144 367334 281232
rect 367442 281144 367622 281232
rect 367730 281144 367910 281232
rect 243214 280928 243394 281016
rect 243502 280928 243682 281016
rect 243790 280928 243970 281016
rect 244078 280928 244258 281016
rect 244366 280928 244546 281016
rect 244654 280928 244834 281016
rect 244942 280928 245122 281016
rect 245230 280928 245410 281016
rect 245664 280928 245844 281016
rect 245952 280928 246132 281016
rect 246240 280928 246420 281016
rect 246528 280928 246708 281016
rect 246816 280928 246996 281016
rect 247104 280928 247284 281016
rect 247392 280928 247572 281016
rect 247680 280928 247860 281016
rect 248114 280928 248294 281016
rect 248402 280928 248582 281016
rect 248690 280928 248870 281016
rect 248978 280928 249158 281016
rect 249266 280928 249446 281016
rect 249554 280928 249734 281016
rect 249842 280928 250022 281016
rect 250130 280928 250310 281016
rect 250564 280928 250744 281016
rect 360436 280928 360560 281016
rect 360814 280928 360994 281016
rect 361102 280928 361282 281016
rect 361390 280928 361570 281016
rect 361678 280928 361858 281016
rect 361966 280928 362146 281016
rect 362254 280928 362434 281016
rect 362542 280928 362722 281016
rect 362830 280928 363010 281016
rect 363264 280928 363444 281016
rect 363552 280928 363732 281016
rect 363840 280928 364020 281016
rect 364128 280928 364308 281016
rect 364416 280928 364596 281016
rect 364704 280928 364884 281016
rect 364992 280928 365172 281016
rect 365280 280928 365460 281016
rect 365714 280928 365894 281016
rect 366002 280928 366182 281016
rect 366290 280928 366470 281016
rect 366578 280928 366758 281016
rect 366866 280928 367046 281016
rect 367154 280928 367334 281016
rect 367442 280928 367622 281016
rect 367730 280928 367910 281016
rect 243214 280452 243394 280540
rect 243502 280452 243682 280540
rect 243790 280452 243970 280540
rect 244078 280452 244258 280540
rect 244366 280452 244546 280540
rect 244654 280452 244834 280540
rect 244942 280452 245122 280540
rect 245230 280452 245410 280540
rect 245664 280452 245844 280540
rect 245952 280452 246132 280540
rect 246240 280452 246420 280540
rect 246528 280452 246708 280540
rect 246816 280452 246996 280540
rect 247104 280452 247284 280540
rect 247392 280452 247572 280540
rect 247680 280452 247860 280540
rect 248114 280452 248294 280540
rect 248402 280452 248582 280540
rect 248690 280452 248870 280540
rect 248978 280452 249158 280540
rect 249266 280452 249446 280540
rect 249554 280452 249734 280540
rect 249842 280452 250022 280540
rect 250130 280452 250310 280540
rect 250564 280452 250744 280540
rect 360436 280452 360560 280540
rect 360814 280452 360994 280540
rect 361102 280452 361282 280540
rect 361390 280452 361570 280540
rect 361678 280452 361858 280540
rect 361966 280452 362146 280540
rect 362254 280452 362434 280540
rect 362542 280452 362722 280540
rect 362830 280452 363010 280540
rect 363264 280452 363444 280540
rect 363552 280452 363732 280540
rect 363840 280452 364020 280540
rect 364128 280452 364308 280540
rect 364416 280452 364596 280540
rect 364704 280452 364884 280540
rect 364992 280452 365172 280540
rect 365280 280452 365460 280540
rect 365714 280452 365894 280540
rect 366002 280452 366182 280540
rect 366290 280452 366470 280540
rect 366578 280452 366758 280540
rect 366866 280452 367046 280540
rect 367154 280452 367334 280540
rect 367442 280452 367622 280540
rect 367730 280452 367910 280540
rect 243214 280236 243394 280324
rect 243502 280236 243682 280324
rect 243790 280236 243970 280324
rect 244078 280236 244258 280324
rect 244366 280236 244546 280324
rect 244654 280236 244834 280324
rect 244942 280236 245122 280324
rect 245230 280236 245410 280324
rect 245664 280236 245844 280324
rect 245952 280236 246132 280324
rect 246240 280236 246420 280324
rect 246528 280236 246708 280324
rect 246816 280236 246996 280324
rect 247104 280236 247284 280324
rect 247392 280236 247572 280324
rect 247680 280236 247860 280324
rect 248114 280236 248294 280324
rect 248402 280236 248582 280324
rect 248690 280236 248870 280324
rect 248978 280236 249158 280324
rect 249266 280236 249446 280324
rect 249554 280236 249734 280324
rect 249842 280236 250022 280324
rect 250130 280236 250310 280324
rect 250564 280236 250744 280324
rect 360436 280236 360560 280324
rect 360814 280236 360994 280324
rect 361102 280236 361282 280324
rect 361390 280236 361570 280324
rect 361678 280236 361858 280324
rect 361966 280236 362146 280324
rect 362254 280236 362434 280324
rect 362542 280236 362722 280324
rect 362830 280236 363010 280324
rect 363264 280236 363444 280324
rect 363552 280236 363732 280324
rect 363840 280236 364020 280324
rect 364128 280236 364308 280324
rect 364416 280236 364596 280324
rect 364704 280236 364884 280324
rect 364992 280236 365172 280324
rect 365280 280236 365460 280324
rect 365714 280236 365894 280324
rect 366002 280236 366182 280324
rect 366290 280236 366470 280324
rect 366578 280236 366758 280324
rect 366866 280236 367046 280324
rect 367154 280236 367334 280324
rect 367442 280236 367622 280324
rect 367730 280236 367910 280324
rect 243214 279760 243394 279848
rect 243502 279760 243682 279848
rect 243790 279760 243970 279848
rect 244078 279760 244258 279848
rect 244366 279760 244546 279848
rect 244654 279760 244834 279848
rect 244942 279760 245122 279848
rect 245230 279760 245410 279848
rect 245664 279760 245844 279848
rect 245952 279760 246132 279848
rect 246240 279760 246420 279848
rect 246528 279760 246708 279848
rect 246816 279760 246996 279848
rect 247104 279760 247284 279848
rect 247392 279760 247572 279848
rect 247680 279760 247860 279848
rect 248114 279760 248294 279848
rect 248402 279760 248582 279848
rect 248690 279760 248870 279848
rect 248978 279760 249158 279848
rect 249266 279760 249446 279848
rect 249554 279760 249734 279848
rect 249842 279760 250022 279848
rect 250130 279760 250310 279848
rect 250564 279760 250744 279848
rect 360436 279760 360560 279848
rect 360814 279760 360994 279848
rect 361102 279760 361282 279848
rect 361390 279760 361570 279848
rect 361678 279760 361858 279848
rect 361966 279760 362146 279848
rect 362254 279760 362434 279848
rect 362542 279760 362722 279848
rect 362830 279760 363010 279848
rect 363264 279760 363444 279848
rect 363552 279760 363732 279848
rect 363840 279760 364020 279848
rect 364128 279760 364308 279848
rect 364416 279760 364596 279848
rect 364704 279760 364884 279848
rect 364992 279760 365172 279848
rect 365280 279760 365460 279848
rect 365714 279760 365894 279848
rect 366002 279760 366182 279848
rect 366290 279760 366470 279848
rect 366578 279760 366758 279848
rect 366866 279760 367046 279848
rect 367154 279760 367334 279848
rect 367442 279760 367622 279848
rect 367730 279760 367910 279848
rect 243214 279544 243394 279632
rect 243502 279544 243682 279632
rect 243790 279544 243970 279632
rect 244078 279544 244258 279632
rect 244366 279544 244546 279632
rect 244654 279544 244834 279632
rect 244942 279544 245122 279632
rect 245230 279544 245410 279632
rect 245664 279544 245844 279632
rect 245952 279544 246132 279632
rect 246240 279544 246420 279632
rect 246528 279544 246708 279632
rect 246816 279544 246996 279632
rect 247104 279544 247284 279632
rect 247392 279544 247572 279632
rect 247680 279544 247860 279632
rect 248114 279544 248294 279632
rect 248402 279544 248582 279632
rect 248690 279544 248870 279632
rect 248978 279544 249158 279632
rect 249266 279544 249446 279632
rect 249554 279544 249734 279632
rect 249842 279544 250022 279632
rect 250130 279544 250310 279632
rect 250564 279544 250744 279632
rect 360436 279544 360560 279632
rect 360814 279544 360994 279632
rect 361102 279544 361282 279632
rect 361390 279544 361570 279632
rect 361678 279544 361858 279632
rect 361966 279544 362146 279632
rect 362254 279544 362434 279632
rect 362542 279544 362722 279632
rect 362830 279544 363010 279632
rect 363264 279544 363444 279632
rect 363552 279544 363732 279632
rect 363840 279544 364020 279632
rect 364128 279544 364308 279632
rect 364416 279544 364596 279632
rect 364704 279544 364884 279632
rect 364992 279544 365172 279632
rect 365280 279544 365460 279632
rect 365714 279544 365894 279632
rect 366002 279544 366182 279632
rect 366290 279544 366470 279632
rect 366578 279544 366758 279632
rect 366866 279544 367046 279632
rect 367154 279544 367334 279632
rect 367442 279544 367622 279632
rect 367730 279544 367910 279632
rect 243214 279068 243394 279156
rect 243502 279068 243682 279156
rect 243790 279068 243970 279156
rect 244078 279068 244258 279156
rect 244366 279068 244546 279156
rect 244654 279068 244834 279156
rect 244942 279068 245122 279156
rect 245230 279068 245410 279156
rect 245664 279068 245844 279156
rect 245952 279068 246132 279156
rect 246240 279068 246420 279156
rect 246528 279068 246708 279156
rect 246816 279068 246996 279156
rect 247104 279068 247284 279156
rect 247392 279068 247572 279156
rect 247680 279068 247860 279156
rect 248114 279068 248294 279156
rect 248402 279068 248582 279156
rect 248690 279068 248870 279156
rect 248978 279068 249158 279156
rect 249266 279068 249446 279156
rect 249554 279068 249734 279156
rect 249842 279068 250022 279156
rect 250130 279068 250310 279156
rect 250564 279068 250744 279156
rect 360436 279068 360560 279156
rect 360814 279068 360994 279156
rect 361102 279068 361282 279156
rect 361390 279068 361570 279156
rect 361678 279068 361858 279156
rect 361966 279068 362146 279156
rect 362254 279068 362434 279156
rect 362542 279068 362722 279156
rect 362830 279068 363010 279156
rect 363264 279068 363444 279156
rect 363552 279068 363732 279156
rect 363840 279068 364020 279156
rect 364128 279068 364308 279156
rect 364416 279068 364596 279156
rect 364704 279068 364884 279156
rect 364992 279068 365172 279156
rect 365280 279068 365460 279156
rect 365714 279068 365894 279156
rect 366002 279068 366182 279156
rect 366290 279068 366470 279156
rect 366578 279068 366758 279156
rect 366866 279068 367046 279156
rect 367154 279068 367334 279156
rect 367442 279068 367622 279156
rect 367730 279068 367910 279156
rect 243214 278594 243394 278682
rect 243502 278594 243682 278682
rect 243790 278594 243970 278682
rect 244078 278594 244258 278682
rect 244366 278594 244546 278682
rect 244654 278594 244834 278682
rect 244942 278594 245122 278682
rect 245230 278594 245410 278682
rect 245664 278594 245844 278682
rect 245952 278594 246132 278682
rect 246240 278594 246420 278682
rect 246528 278594 246708 278682
rect 246816 278594 246996 278682
rect 247104 278594 247284 278682
rect 247392 278594 247572 278682
rect 247680 278594 247860 278682
rect 248114 278594 248294 278682
rect 248402 278594 248582 278682
rect 248690 278594 248870 278682
rect 248978 278594 249158 278682
rect 249266 278594 249446 278682
rect 249554 278594 249734 278682
rect 249842 278594 250022 278682
rect 250130 278594 250310 278682
rect 250564 278594 250744 278682
rect 360436 278594 360560 278682
rect 360814 278594 360994 278682
rect 361102 278594 361282 278682
rect 361390 278594 361570 278682
rect 361678 278594 361858 278682
rect 361966 278594 362146 278682
rect 362254 278594 362434 278682
rect 362542 278594 362722 278682
rect 362830 278594 363010 278682
rect 363264 278594 363444 278682
rect 363552 278594 363732 278682
rect 363840 278594 364020 278682
rect 364128 278594 364308 278682
rect 364416 278594 364596 278682
rect 364704 278594 364884 278682
rect 364992 278594 365172 278682
rect 365280 278594 365460 278682
rect 365714 278594 365894 278682
rect 366002 278594 366182 278682
rect 366290 278594 366470 278682
rect 366578 278594 366758 278682
rect 366866 278594 367046 278682
rect 367154 278594 367334 278682
rect 367442 278594 367622 278682
rect 367730 278594 367910 278682
rect 243214 278118 243394 278206
rect 243502 278118 243682 278206
rect 243790 278118 243970 278206
rect 244078 278118 244258 278206
rect 244366 278118 244546 278206
rect 244654 278118 244834 278206
rect 244942 278118 245122 278206
rect 245230 278118 245410 278206
rect 245664 278118 245844 278206
rect 245952 278118 246132 278206
rect 246240 278118 246420 278206
rect 246528 278118 246708 278206
rect 246816 278118 246996 278206
rect 247104 278118 247284 278206
rect 247392 278118 247572 278206
rect 247680 278118 247860 278206
rect 248114 278118 248294 278206
rect 248402 278118 248582 278206
rect 248690 278118 248870 278206
rect 248978 278118 249158 278206
rect 249266 278118 249446 278206
rect 249554 278118 249734 278206
rect 249842 278118 250022 278206
rect 250130 278118 250310 278206
rect 250564 278118 250744 278206
rect 360436 278118 360560 278206
rect 360814 278118 360994 278206
rect 361102 278118 361282 278206
rect 361390 278118 361570 278206
rect 361678 278118 361858 278206
rect 361966 278118 362146 278206
rect 362254 278118 362434 278206
rect 362542 278118 362722 278206
rect 362830 278118 363010 278206
rect 363264 278118 363444 278206
rect 363552 278118 363732 278206
rect 363840 278118 364020 278206
rect 364128 278118 364308 278206
rect 364416 278118 364596 278206
rect 364704 278118 364884 278206
rect 364992 278118 365172 278206
rect 365280 278118 365460 278206
rect 365714 278118 365894 278206
rect 366002 278118 366182 278206
rect 366290 278118 366470 278206
rect 366578 278118 366758 278206
rect 366866 278118 367046 278206
rect 367154 278118 367334 278206
rect 367442 278118 367622 278206
rect 367730 278118 367910 278206
rect 243214 277902 243394 277990
rect 243502 277902 243682 277990
rect 243790 277902 243970 277990
rect 244078 277902 244258 277990
rect 244366 277902 244546 277990
rect 244654 277902 244834 277990
rect 244942 277902 245122 277990
rect 245230 277902 245410 277990
rect 245664 277902 245844 277990
rect 245952 277902 246132 277990
rect 246240 277902 246420 277990
rect 246528 277902 246708 277990
rect 246816 277902 246996 277990
rect 247104 277902 247284 277990
rect 247392 277902 247572 277990
rect 247680 277902 247860 277990
rect 248114 277902 248294 277990
rect 248402 277902 248582 277990
rect 248690 277902 248870 277990
rect 248978 277902 249158 277990
rect 249266 277902 249446 277990
rect 249554 277902 249734 277990
rect 249842 277902 250022 277990
rect 250130 277902 250310 277990
rect 250564 277902 250744 277990
rect 360436 277902 360560 277990
rect 360814 277902 360994 277990
rect 361102 277902 361282 277990
rect 361390 277902 361570 277990
rect 361678 277902 361858 277990
rect 361966 277902 362146 277990
rect 362254 277902 362434 277990
rect 362542 277902 362722 277990
rect 362830 277902 363010 277990
rect 363264 277902 363444 277990
rect 363552 277902 363732 277990
rect 363840 277902 364020 277990
rect 364128 277902 364308 277990
rect 364416 277902 364596 277990
rect 364704 277902 364884 277990
rect 364992 277902 365172 277990
rect 365280 277902 365460 277990
rect 365714 277902 365894 277990
rect 366002 277902 366182 277990
rect 366290 277902 366470 277990
rect 366578 277902 366758 277990
rect 366866 277902 367046 277990
rect 367154 277902 367334 277990
rect 367442 277902 367622 277990
rect 367730 277902 367910 277990
rect 243214 277426 243394 277514
rect 243502 277426 243682 277514
rect 243790 277426 243970 277514
rect 244078 277426 244258 277514
rect 244366 277426 244546 277514
rect 244654 277426 244834 277514
rect 244942 277426 245122 277514
rect 245230 277426 245410 277514
rect 245664 277426 245844 277514
rect 245952 277426 246132 277514
rect 246240 277426 246420 277514
rect 246528 277426 246708 277514
rect 246816 277426 246996 277514
rect 247104 277426 247284 277514
rect 247392 277426 247572 277514
rect 247680 277426 247860 277514
rect 248114 277426 248294 277514
rect 248402 277426 248582 277514
rect 248690 277426 248870 277514
rect 248978 277426 249158 277514
rect 249266 277426 249446 277514
rect 249554 277426 249734 277514
rect 249842 277426 250022 277514
rect 250130 277426 250310 277514
rect 250564 277426 250744 277514
rect 360436 277426 360560 277514
rect 360814 277426 360994 277514
rect 361102 277426 361282 277514
rect 361390 277426 361570 277514
rect 361678 277426 361858 277514
rect 361966 277426 362146 277514
rect 362254 277426 362434 277514
rect 362542 277426 362722 277514
rect 362830 277426 363010 277514
rect 363264 277426 363444 277514
rect 363552 277426 363732 277514
rect 363840 277426 364020 277514
rect 364128 277426 364308 277514
rect 364416 277426 364596 277514
rect 364704 277426 364884 277514
rect 364992 277426 365172 277514
rect 365280 277426 365460 277514
rect 365714 277426 365894 277514
rect 366002 277426 366182 277514
rect 366290 277426 366470 277514
rect 366578 277426 366758 277514
rect 366866 277426 367046 277514
rect 367154 277426 367334 277514
rect 367442 277426 367622 277514
rect 367730 277426 367910 277514
rect 243214 277210 243394 277298
rect 243502 277210 243682 277298
rect 243790 277210 243970 277298
rect 244078 277210 244258 277298
rect 244366 277210 244546 277298
rect 244654 277210 244834 277298
rect 244942 277210 245122 277298
rect 245230 277210 245410 277298
rect 245664 277210 245844 277298
rect 245952 277210 246132 277298
rect 246240 277210 246420 277298
rect 246528 277210 246708 277298
rect 246816 277210 246996 277298
rect 247104 277210 247284 277298
rect 247392 277210 247572 277298
rect 247680 277210 247860 277298
rect 248114 277210 248294 277298
rect 248402 277210 248582 277298
rect 248690 277210 248870 277298
rect 248978 277210 249158 277298
rect 249266 277210 249446 277298
rect 249554 277210 249734 277298
rect 249842 277210 250022 277298
rect 250130 277210 250310 277298
rect 250564 277210 250744 277298
rect 360436 277210 360560 277298
rect 360814 277210 360994 277298
rect 361102 277210 361282 277298
rect 361390 277210 361570 277298
rect 361678 277210 361858 277298
rect 361966 277210 362146 277298
rect 362254 277210 362434 277298
rect 362542 277210 362722 277298
rect 362830 277210 363010 277298
rect 363264 277210 363444 277298
rect 363552 277210 363732 277298
rect 363840 277210 364020 277298
rect 364128 277210 364308 277298
rect 364416 277210 364596 277298
rect 364704 277210 364884 277298
rect 364992 277210 365172 277298
rect 365280 277210 365460 277298
rect 365714 277210 365894 277298
rect 366002 277210 366182 277298
rect 366290 277210 366470 277298
rect 366578 277210 366758 277298
rect 366866 277210 367046 277298
rect 367154 277210 367334 277298
rect 367442 277210 367622 277298
rect 367730 277210 367910 277298
rect 243214 276734 243394 276822
rect 243502 276734 243682 276822
rect 243790 276734 243970 276822
rect 244078 276734 244258 276822
rect 244366 276734 244546 276822
rect 244654 276734 244834 276822
rect 244942 276734 245122 276822
rect 245230 276734 245410 276822
rect 245664 276734 245844 276822
rect 245952 276734 246132 276822
rect 246240 276734 246420 276822
rect 246528 276734 246708 276822
rect 246816 276734 246996 276822
rect 247104 276734 247284 276822
rect 247392 276734 247572 276822
rect 247680 276734 247860 276822
rect 248114 276734 248294 276822
rect 248402 276734 248582 276822
rect 248690 276734 248870 276822
rect 248978 276734 249158 276822
rect 249266 276734 249446 276822
rect 249554 276734 249734 276822
rect 249842 276734 250022 276822
rect 250130 276734 250310 276822
rect 250564 276734 250744 276822
rect 360436 276734 360560 276822
rect 360814 276734 360994 276822
rect 361102 276734 361282 276822
rect 361390 276734 361570 276822
rect 361678 276734 361858 276822
rect 361966 276734 362146 276822
rect 362254 276734 362434 276822
rect 362542 276734 362722 276822
rect 362830 276734 363010 276822
rect 363264 276734 363444 276822
rect 363552 276734 363732 276822
rect 363840 276734 364020 276822
rect 364128 276734 364308 276822
rect 364416 276734 364596 276822
rect 364704 276734 364884 276822
rect 364992 276734 365172 276822
rect 365280 276734 365460 276822
rect 365714 276734 365894 276822
rect 366002 276734 366182 276822
rect 366290 276734 366470 276822
rect 366578 276734 366758 276822
rect 366866 276734 367046 276822
rect 367154 276734 367334 276822
rect 367442 276734 367622 276822
rect 367730 276734 367910 276822
rect 243214 276518 243394 276606
rect 243502 276518 243682 276606
rect 243790 276518 243970 276606
rect 244078 276518 244258 276606
rect 244366 276518 244546 276606
rect 244654 276518 244834 276606
rect 244942 276518 245122 276606
rect 245230 276518 245410 276606
rect 245664 276518 245844 276606
rect 245952 276518 246132 276606
rect 246240 276518 246420 276606
rect 246528 276518 246708 276606
rect 246816 276518 246996 276606
rect 247104 276518 247284 276606
rect 247392 276518 247572 276606
rect 247680 276518 247860 276606
rect 248114 276518 248294 276606
rect 248402 276518 248582 276606
rect 248690 276518 248870 276606
rect 248978 276518 249158 276606
rect 249266 276518 249446 276606
rect 249554 276518 249734 276606
rect 249842 276518 250022 276606
rect 250130 276518 250310 276606
rect 250564 276518 250744 276606
rect 360436 276518 360560 276606
rect 360814 276518 360994 276606
rect 361102 276518 361282 276606
rect 361390 276518 361570 276606
rect 361678 276518 361858 276606
rect 361966 276518 362146 276606
rect 362254 276518 362434 276606
rect 362542 276518 362722 276606
rect 362830 276518 363010 276606
rect 363264 276518 363444 276606
rect 363552 276518 363732 276606
rect 363840 276518 364020 276606
rect 364128 276518 364308 276606
rect 364416 276518 364596 276606
rect 364704 276518 364884 276606
rect 364992 276518 365172 276606
rect 365280 276518 365460 276606
rect 365714 276518 365894 276606
rect 366002 276518 366182 276606
rect 366290 276518 366470 276606
rect 366578 276518 366758 276606
rect 366866 276518 367046 276606
rect 367154 276518 367334 276606
rect 367442 276518 367622 276606
rect 367730 276518 367910 276606
rect 243214 276042 243394 276130
rect 243502 276042 243682 276130
rect 243790 276042 243970 276130
rect 244078 276042 244258 276130
rect 244366 276042 244546 276130
rect 244654 276042 244834 276130
rect 244942 276042 245122 276130
rect 245230 276042 245410 276130
rect 245664 276042 245844 276130
rect 245952 276042 246132 276130
rect 246240 276042 246420 276130
rect 246528 276042 246708 276130
rect 246816 276042 246996 276130
rect 247104 276042 247284 276130
rect 247392 276042 247572 276130
rect 247680 276042 247860 276130
rect 248114 276042 248294 276130
rect 248402 276042 248582 276130
rect 248690 276042 248870 276130
rect 248978 276042 249158 276130
rect 249266 276042 249446 276130
rect 249554 276042 249734 276130
rect 249842 276042 250022 276130
rect 250130 276042 250310 276130
rect 250564 276042 250744 276130
rect 360436 276042 360560 276130
rect 360814 276042 360994 276130
rect 361102 276042 361282 276130
rect 361390 276042 361570 276130
rect 361678 276042 361858 276130
rect 361966 276042 362146 276130
rect 362254 276042 362434 276130
rect 362542 276042 362722 276130
rect 362830 276042 363010 276130
rect 363264 276042 363444 276130
rect 363552 276042 363732 276130
rect 363840 276042 364020 276130
rect 364128 276042 364308 276130
rect 364416 276042 364596 276130
rect 364704 276042 364884 276130
rect 364992 276042 365172 276130
rect 365280 276042 365460 276130
rect 365714 276042 365894 276130
rect 366002 276042 366182 276130
rect 366290 276042 366470 276130
rect 366578 276042 366758 276130
rect 366866 276042 367046 276130
rect 367154 276042 367334 276130
rect 367442 276042 367622 276130
rect 367730 276042 367910 276130
rect 243214 275568 243394 275656
rect 243502 275568 243682 275656
rect 243790 275568 243970 275656
rect 244078 275568 244258 275656
rect 244366 275568 244546 275656
rect 244654 275568 244834 275656
rect 244942 275568 245122 275656
rect 245230 275568 245410 275656
rect 245664 275568 245844 275656
rect 245952 275568 246132 275656
rect 246240 275568 246420 275656
rect 246528 275568 246708 275656
rect 246816 275568 246996 275656
rect 247104 275568 247284 275656
rect 247392 275568 247572 275656
rect 247680 275568 247860 275656
rect 248114 275568 248294 275656
rect 248402 275568 248582 275656
rect 248690 275568 248870 275656
rect 248978 275568 249158 275656
rect 249266 275568 249446 275656
rect 249554 275568 249734 275656
rect 249842 275568 250022 275656
rect 250130 275568 250310 275656
rect 250564 275568 250744 275656
rect 360436 275568 360560 275656
rect 360814 275568 360994 275656
rect 361102 275568 361282 275656
rect 361390 275568 361570 275656
rect 361678 275568 361858 275656
rect 361966 275568 362146 275656
rect 362254 275568 362434 275656
rect 362542 275568 362722 275656
rect 362830 275568 363010 275656
rect 363264 275568 363444 275656
rect 363552 275568 363732 275656
rect 363840 275568 364020 275656
rect 364128 275568 364308 275656
rect 364416 275568 364596 275656
rect 364704 275568 364884 275656
rect 364992 275568 365172 275656
rect 365280 275568 365460 275656
rect 365714 275568 365894 275656
rect 366002 275568 366182 275656
rect 366290 275568 366470 275656
rect 366578 275568 366758 275656
rect 366866 275568 367046 275656
rect 367154 275568 367334 275656
rect 367442 275568 367622 275656
rect 367730 275568 367910 275656
rect 243214 275092 243394 275180
rect 243502 275092 243682 275180
rect 243790 275092 243970 275180
rect 244078 275092 244258 275180
rect 244366 275092 244546 275180
rect 244654 275092 244834 275180
rect 244942 275092 245122 275180
rect 245230 275092 245410 275180
rect 245664 275092 245844 275180
rect 245952 275092 246132 275180
rect 246240 275092 246420 275180
rect 246528 275092 246708 275180
rect 246816 275092 246996 275180
rect 247104 275092 247284 275180
rect 247392 275092 247572 275180
rect 247680 275092 247860 275180
rect 248114 275092 248294 275180
rect 248402 275092 248582 275180
rect 248690 275092 248870 275180
rect 248978 275092 249158 275180
rect 249266 275092 249446 275180
rect 249554 275092 249734 275180
rect 249842 275092 250022 275180
rect 250130 275092 250310 275180
rect 250564 275092 250744 275180
rect 360436 275092 360560 275180
rect 360814 275092 360994 275180
rect 361102 275092 361282 275180
rect 361390 275092 361570 275180
rect 361678 275092 361858 275180
rect 361966 275092 362146 275180
rect 362254 275092 362434 275180
rect 362542 275092 362722 275180
rect 362830 275092 363010 275180
rect 363264 275092 363444 275180
rect 363552 275092 363732 275180
rect 363840 275092 364020 275180
rect 364128 275092 364308 275180
rect 364416 275092 364596 275180
rect 364704 275092 364884 275180
rect 364992 275092 365172 275180
rect 365280 275092 365460 275180
rect 365714 275092 365894 275180
rect 366002 275092 366182 275180
rect 366290 275092 366470 275180
rect 366578 275092 366758 275180
rect 366866 275092 367046 275180
rect 367154 275092 367334 275180
rect 367442 275092 367622 275180
rect 367730 275092 367910 275180
rect 243214 274876 243394 274964
rect 243502 274876 243682 274964
rect 243790 274876 243970 274964
rect 244078 274876 244258 274964
rect 244366 274876 244546 274964
rect 244654 274876 244834 274964
rect 244942 274876 245122 274964
rect 245230 274876 245410 274964
rect 245664 274876 245844 274964
rect 245952 274876 246132 274964
rect 246240 274876 246420 274964
rect 246528 274876 246708 274964
rect 246816 274876 246996 274964
rect 247104 274876 247284 274964
rect 247392 274876 247572 274964
rect 247680 274876 247860 274964
rect 248114 274876 248294 274964
rect 248402 274876 248582 274964
rect 248690 274876 248870 274964
rect 248978 274876 249158 274964
rect 249266 274876 249446 274964
rect 249554 274876 249734 274964
rect 249842 274876 250022 274964
rect 250130 274876 250310 274964
rect 250564 274876 250744 274964
rect 360436 274876 360560 274964
rect 360814 274876 360994 274964
rect 361102 274876 361282 274964
rect 361390 274876 361570 274964
rect 361678 274876 361858 274964
rect 361966 274876 362146 274964
rect 362254 274876 362434 274964
rect 362542 274876 362722 274964
rect 362830 274876 363010 274964
rect 363264 274876 363444 274964
rect 363552 274876 363732 274964
rect 363840 274876 364020 274964
rect 364128 274876 364308 274964
rect 364416 274876 364596 274964
rect 364704 274876 364884 274964
rect 364992 274876 365172 274964
rect 365280 274876 365460 274964
rect 365714 274876 365894 274964
rect 366002 274876 366182 274964
rect 366290 274876 366470 274964
rect 366578 274876 366758 274964
rect 366866 274876 367046 274964
rect 367154 274876 367334 274964
rect 367442 274876 367622 274964
rect 367730 274876 367910 274964
rect 243214 274400 243394 274488
rect 243502 274400 243682 274488
rect 243790 274400 243970 274488
rect 244078 274400 244258 274488
rect 244366 274400 244546 274488
rect 244654 274400 244834 274488
rect 244942 274400 245122 274488
rect 245230 274400 245410 274488
rect 245664 274400 245844 274488
rect 245952 274400 246132 274488
rect 246240 274400 246420 274488
rect 246528 274400 246708 274488
rect 246816 274400 246996 274488
rect 247104 274400 247284 274488
rect 247392 274400 247572 274488
rect 247680 274400 247860 274488
rect 248114 274400 248294 274488
rect 248402 274400 248582 274488
rect 248690 274400 248870 274488
rect 248978 274400 249158 274488
rect 249266 274400 249446 274488
rect 249554 274400 249734 274488
rect 249842 274400 250022 274488
rect 250130 274400 250310 274488
rect 250564 274400 250744 274488
rect 360436 274400 360560 274488
rect 360814 274400 360994 274488
rect 361102 274400 361282 274488
rect 361390 274400 361570 274488
rect 361678 274400 361858 274488
rect 361966 274400 362146 274488
rect 362254 274400 362434 274488
rect 362542 274400 362722 274488
rect 362830 274400 363010 274488
rect 363264 274400 363444 274488
rect 363552 274400 363732 274488
rect 363840 274400 364020 274488
rect 364128 274400 364308 274488
rect 364416 274400 364596 274488
rect 364704 274400 364884 274488
rect 364992 274400 365172 274488
rect 365280 274400 365460 274488
rect 365714 274400 365894 274488
rect 366002 274400 366182 274488
rect 366290 274400 366470 274488
rect 366578 274400 366758 274488
rect 366866 274400 367046 274488
rect 367154 274400 367334 274488
rect 367442 274400 367622 274488
rect 367730 274400 367910 274488
rect 243214 274184 243394 274272
rect 243502 274184 243682 274272
rect 243790 274184 243970 274272
rect 244078 274184 244258 274272
rect 244366 274184 244546 274272
rect 244654 274184 244834 274272
rect 244942 274184 245122 274272
rect 245230 274184 245410 274272
rect 245664 274184 245844 274272
rect 245952 274184 246132 274272
rect 246240 274184 246420 274272
rect 246528 274184 246708 274272
rect 246816 274184 246996 274272
rect 247104 274184 247284 274272
rect 247392 274184 247572 274272
rect 247680 274184 247860 274272
rect 248114 274184 248294 274272
rect 248402 274184 248582 274272
rect 248690 274184 248870 274272
rect 248978 274184 249158 274272
rect 249266 274184 249446 274272
rect 249554 274184 249734 274272
rect 249842 274184 250022 274272
rect 250130 274184 250310 274272
rect 250564 274184 250744 274272
rect 360436 274184 360560 274272
rect 360814 274184 360994 274272
rect 361102 274184 361282 274272
rect 361390 274184 361570 274272
rect 361678 274184 361858 274272
rect 361966 274184 362146 274272
rect 362254 274184 362434 274272
rect 362542 274184 362722 274272
rect 362830 274184 363010 274272
rect 363264 274184 363444 274272
rect 363552 274184 363732 274272
rect 363840 274184 364020 274272
rect 364128 274184 364308 274272
rect 364416 274184 364596 274272
rect 364704 274184 364884 274272
rect 364992 274184 365172 274272
rect 365280 274184 365460 274272
rect 365714 274184 365894 274272
rect 366002 274184 366182 274272
rect 366290 274184 366470 274272
rect 366578 274184 366758 274272
rect 366866 274184 367046 274272
rect 367154 274184 367334 274272
rect 367442 274184 367622 274272
rect 367730 274184 367910 274272
rect 243214 273708 243394 273796
rect 243502 273708 243682 273796
rect 243790 273708 243970 273796
rect 244078 273708 244258 273796
rect 244366 273708 244546 273796
rect 244654 273708 244834 273796
rect 244942 273708 245122 273796
rect 245230 273708 245410 273796
rect 245664 273708 245844 273796
rect 245952 273708 246132 273796
rect 246240 273708 246420 273796
rect 246528 273708 246708 273796
rect 246816 273708 246996 273796
rect 247104 273708 247284 273796
rect 247392 273708 247572 273796
rect 247680 273708 247860 273796
rect 248114 273708 248294 273796
rect 248402 273708 248582 273796
rect 248690 273708 248870 273796
rect 248978 273708 249158 273796
rect 249266 273708 249446 273796
rect 249554 273708 249734 273796
rect 249842 273708 250022 273796
rect 250130 273708 250310 273796
rect 250564 273708 250744 273796
rect 360436 273708 360560 273796
rect 360814 273708 360994 273796
rect 361102 273708 361282 273796
rect 361390 273708 361570 273796
rect 361678 273708 361858 273796
rect 361966 273708 362146 273796
rect 362254 273708 362434 273796
rect 362542 273708 362722 273796
rect 362830 273708 363010 273796
rect 363264 273708 363444 273796
rect 363552 273708 363732 273796
rect 363840 273708 364020 273796
rect 364128 273708 364308 273796
rect 364416 273708 364596 273796
rect 364704 273708 364884 273796
rect 364992 273708 365172 273796
rect 365280 273708 365460 273796
rect 365714 273708 365894 273796
rect 366002 273708 366182 273796
rect 366290 273708 366470 273796
rect 366578 273708 366758 273796
rect 366866 273708 367046 273796
rect 367154 273708 367334 273796
rect 367442 273708 367622 273796
rect 367730 273708 367910 273796
rect 243214 273492 243394 273580
rect 243502 273492 243682 273580
rect 243790 273492 243970 273580
rect 244078 273492 244258 273580
rect 244366 273492 244546 273580
rect 244654 273492 244834 273580
rect 244942 273492 245122 273580
rect 245230 273492 245410 273580
rect 245664 273492 245844 273580
rect 245952 273492 246132 273580
rect 246240 273492 246420 273580
rect 246528 273492 246708 273580
rect 246816 273492 246996 273580
rect 247104 273492 247284 273580
rect 247392 273492 247572 273580
rect 247680 273492 247860 273580
rect 248114 273492 248294 273580
rect 248402 273492 248582 273580
rect 248690 273492 248870 273580
rect 248978 273492 249158 273580
rect 249266 273492 249446 273580
rect 249554 273492 249734 273580
rect 249842 273492 250022 273580
rect 250130 273492 250310 273580
rect 250564 273492 250744 273580
rect 360436 273492 360560 273580
rect 360814 273492 360994 273580
rect 361102 273492 361282 273580
rect 361390 273492 361570 273580
rect 361678 273492 361858 273580
rect 361966 273492 362146 273580
rect 362254 273492 362434 273580
rect 362542 273492 362722 273580
rect 362830 273492 363010 273580
rect 363264 273492 363444 273580
rect 363552 273492 363732 273580
rect 363840 273492 364020 273580
rect 364128 273492 364308 273580
rect 364416 273492 364596 273580
rect 364704 273492 364884 273580
rect 364992 273492 365172 273580
rect 365280 273492 365460 273580
rect 365714 273492 365894 273580
rect 366002 273492 366182 273580
rect 366290 273492 366470 273580
rect 366578 273492 366758 273580
rect 366866 273492 367046 273580
rect 367154 273492 367334 273580
rect 367442 273492 367622 273580
rect 367730 273492 367910 273580
rect 243214 273016 243394 273104
rect 243502 273016 243682 273104
rect 243790 273016 243970 273104
rect 244078 273016 244258 273104
rect 244366 273016 244546 273104
rect 244654 273016 244834 273104
rect 244942 273016 245122 273104
rect 245230 273016 245410 273104
rect 245664 273016 245844 273104
rect 245952 273016 246132 273104
rect 246240 273016 246420 273104
rect 246528 273016 246708 273104
rect 246816 273016 246996 273104
rect 247104 273016 247284 273104
rect 247392 273016 247572 273104
rect 247680 273016 247860 273104
rect 248114 273016 248294 273104
rect 248402 273016 248582 273104
rect 248690 273016 248870 273104
rect 248978 273016 249158 273104
rect 249266 273016 249446 273104
rect 249554 273016 249734 273104
rect 249842 273016 250022 273104
rect 250130 273016 250310 273104
rect 250564 273016 250744 273104
rect 360436 273016 360560 273104
rect 360814 273016 360994 273104
rect 361102 273016 361282 273104
rect 361390 273016 361570 273104
rect 361678 273016 361858 273104
rect 361966 273016 362146 273104
rect 362254 273016 362434 273104
rect 362542 273016 362722 273104
rect 362830 273016 363010 273104
rect 363264 273016 363444 273104
rect 363552 273016 363732 273104
rect 363840 273016 364020 273104
rect 364128 273016 364308 273104
rect 364416 273016 364596 273104
rect 364704 273016 364884 273104
rect 364992 273016 365172 273104
rect 365280 273016 365460 273104
rect 365714 273016 365894 273104
rect 366002 273016 366182 273104
rect 366290 273016 366470 273104
rect 366578 273016 366758 273104
rect 366866 273016 367046 273104
rect 367154 273016 367334 273104
rect 367442 273016 367622 273104
rect 367730 273016 367910 273104
rect 243214 272542 243394 272630
rect 243502 272542 243682 272630
rect 243790 272542 243970 272630
rect 244078 272542 244258 272630
rect 244366 272542 244546 272630
rect 244654 272542 244834 272630
rect 244942 272542 245122 272630
rect 245230 272542 245410 272630
rect 245664 272542 245844 272630
rect 245952 272542 246132 272630
rect 246240 272542 246420 272630
rect 246528 272542 246708 272630
rect 246816 272542 246996 272630
rect 247104 272542 247284 272630
rect 247392 272542 247572 272630
rect 247680 272542 247860 272630
rect 248114 272542 248294 272630
rect 248402 272542 248582 272630
rect 248690 272542 248870 272630
rect 248978 272542 249158 272630
rect 249266 272542 249446 272630
rect 249554 272542 249734 272630
rect 249842 272542 250022 272630
rect 250130 272542 250310 272630
rect 250564 272542 250744 272630
rect 360436 272542 360560 272630
rect 360814 272542 360994 272630
rect 361102 272542 361282 272630
rect 361390 272542 361570 272630
rect 361678 272542 361858 272630
rect 361966 272542 362146 272630
rect 362254 272542 362434 272630
rect 362542 272542 362722 272630
rect 362830 272542 363010 272630
rect 363264 272542 363444 272630
rect 363552 272542 363732 272630
rect 363840 272542 364020 272630
rect 364128 272542 364308 272630
rect 364416 272542 364596 272630
rect 364704 272542 364884 272630
rect 364992 272542 365172 272630
rect 365280 272542 365460 272630
rect 365714 272542 365894 272630
rect 366002 272542 366182 272630
rect 366290 272542 366470 272630
rect 366578 272542 366758 272630
rect 366866 272542 367046 272630
rect 367154 272542 367334 272630
rect 367442 272542 367622 272630
rect 367730 272542 367910 272630
rect 243214 272066 243394 272154
rect 243502 272066 243682 272154
rect 243790 272066 243970 272154
rect 244078 272066 244258 272154
rect 244366 272066 244546 272154
rect 244654 272066 244834 272154
rect 244942 272066 245122 272154
rect 245230 272066 245410 272154
rect 245664 272066 245844 272154
rect 245952 272066 246132 272154
rect 246240 272066 246420 272154
rect 246528 272066 246708 272154
rect 246816 272066 246996 272154
rect 247104 272066 247284 272154
rect 247392 272066 247572 272154
rect 247680 272066 247860 272154
rect 248114 272066 248294 272154
rect 248402 272066 248582 272154
rect 248690 272066 248870 272154
rect 248978 272066 249158 272154
rect 249266 272066 249446 272154
rect 249554 272066 249734 272154
rect 249842 272066 250022 272154
rect 250130 272066 250310 272154
rect 250564 272066 250744 272154
rect 360436 272066 360560 272154
rect 360814 272066 360994 272154
rect 361102 272066 361282 272154
rect 361390 272066 361570 272154
rect 361678 272066 361858 272154
rect 361966 272066 362146 272154
rect 362254 272066 362434 272154
rect 362542 272066 362722 272154
rect 362830 272066 363010 272154
rect 363264 272066 363444 272154
rect 363552 272066 363732 272154
rect 363840 272066 364020 272154
rect 364128 272066 364308 272154
rect 364416 272066 364596 272154
rect 364704 272066 364884 272154
rect 364992 272066 365172 272154
rect 365280 272066 365460 272154
rect 365714 272066 365894 272154
rect 366002 272066 366182 272154
rect 366290 272066 366470 272154
rect 366578 272066 366758 272154
rect 366866 272066 367046 272154
rect 367154 272066 367334 272154
rect 367442 272066 367622 272154
rect 367730 272066 367910 272154
rect 243214 271850 243394 271938
rect 243502 271850 243682 271938
rect 243790 271850 243970 271938
rect 244078 271850 244258 271938
rect 244366 271850 244546 271938
rect 244654 271850 244834 271938
rect 244942 271850 245122 271938
rect 245230 271850 245410 271938
rect 245664 271850 245844 271938
rect 245952 271850 246132 271938
rect 246240 271850 246420 271938
rect 246528 271850 246708 271938
rect 246816 271850 246996 271938
rect 247104 271850 247284 271938
rect 247392 271850 247572 271938
rect 247680 271850 247860 271938
rect 248114 271850 248294 271938
rect 248402 271850 248582 271938
rect 248690 271850 248870 271938
rect 248978 271850 249158 271938
rect 249266 271850 249446 271938
rect 249554 271850 249734 271938
rect 249842 271850 250022 271938
rect 250130 271850 250310 271938
rect 250564 271850 250744 271938
rect 360436 271850 360560 271938
rect 360814 271850 360994 271938
rect 361102 271850 361282 271938
rect 361390 271850 361570 271938
rect 361678 271850 361858 271938
rect 361966 271850 362146 271938
rect 362254 271850 362434 271938
rect 362542 271850 362722 271938
rect 362830 271850 363010 271938
rect 363264 271850 363444 271938
rect 363552 271850 363732 271938
rect 363840 271850 364020 271938
rect 364128 271850 364308 271938
rect 364416 271850 364596 271938
rect 364704 271850 364884 271938
rect 364992 271850 365172 271938
rect 365280 271850 365460 271938
rect 365714 271850 365894 271938
rect 366002 271850 366182 271938
rect 366290 271850 366470 271938
rect 366578 271850 366758 271938
rect 366866 271850 367046 271938
rect 367154 271850 367334 271938
rect 367442 271850 367622 271938
rect 367730 271850 367910 271938
rect 243214 271374 243394 271462
rect 243502 271374 243682 271462
rect 243790 271374 243970 271462
rect 244078 271374 244258 271462
rect 244366 271374 244546 271462
rect 244654 271374 244834 271462
rect 244942 271374 245122 271462
rect 245230 271374 245410 271462
rect 245664 271374 245844 271462
rect 245952 271374 246132 271462
rect 246240 271374 246420 271462
rect 246528 271374 246708 271462
rect 246816 271374 246996 271462
rect 247104 271374 247284 271462
rect 247392 271374 247572 271462
rect 247680 271374 247860 271462
rect 248114 271374 248294 271462
rect 248402 271374 248582 271462
rect 248690 271374 248870 271462
rect 248978 271374 249158 271462
rect 249266 271374 249446 271462
rect 249554 271374 249734 271462
rect 249842 271374 250022 271462
rect 250130 271374 250310 271462
rect 250564 271374 250744 271462
rect 360436 271374 360560 271462
rect 360814 271374 360994 271462
rect 361102 271374 361282 271462
rect 361390 271374 361570 271462
rect 361678 271374 361858 271462
rect 361966 271374 362146 271462
rect 362254 271374 362434 271462
rect 362542 271374 362722 271462
rect 362830 271374 363010 271462
rect 363264 271374 363444 271462
rect 363552 271374 363732 271462
rect 363840 271374 364020 271462
rect 364128 271374 364308 271462
rect 364416 271374 364596 271462
rect 364704 271374 364884 271462
rect 364992 271374 365172 271462
rect 365280 271374 365460 271462
rect 365714 271374 365894 271462
rect 366002 271374 366182 271462
rect 366290 271374 366470 271462
rect 366578 271374 366758 271462
rect 366866 271374 367046 271462
rect 367154 271374 367334 271462
rect 367442 271374 367622 271462
rect 367730 271374 367910 271462
rect 243214 271158 243394 271246
rect 243502 271158 243682 271246
rect 243790 271158 243970 271246
rect 244078 271158 244258 271246
rect 244366 271158 244546 271246
rect 244654 271158 244834 271246
rect 244942 271158 245122 271246
rect 245230 271158 245410 271246
rect 245664 271158 245844 271246
rect 245952 271158 246132 271246
rect 246240 271158 246420 271246
rect 246528 271158 246708 271246
rect 246816 271158 246996 271246
rect 247104 271158 247284 271246
rect 247392 271158 247572 271246
rect 247680 271158 247860 271246
rect 248114 271158 248294 271246
rect 248402 271158 248582 271246
rect 248690 271158 248870 271246
rect 248978 271158 249158 271246
rect 249266 271158 249446 271246
rect 249554 271158 249734 271246
rect 249842 271158 250022 271246
rect 250130 271158 250310 271246
rect 250564 271158 250744 271246
rect 360436 271158 360560 271246
rect 360814 271158 360994 271246
rect 361102 271158 361282 271246
rect 361390 271158 361570 271246
rect 361678 271158 361858 271246
rect 361966 271158 362146 271246
rect 362254 271158 362434 271246
rect 362542 271158 362722 271246
rect 362830 271158 363010 271246
rect 363264 271158 363444 271246
rect 363552 271158 363732 271246
rect 363840 271158 364020 271246
rect 364128 271158 364308 271246
rect 364416 271158 364596 271246
rect 364704 271158 364884 271246
rect 364992 271158 365172 271246
rect 365280 271158 365460 271246
rect 365714 271158 365894 271246
rect 366002 271158 366182 271246
rect 366290 271158 366470 271246
rect 366578 271158 366758 271246
rect 366866 271158 367046 271246
rect 367154 271158 367334 271246
rect 367442 271158 367622 271246
rect 367730 271158 367910 271246
rect 243214 270682 243394 270770
rect 243502 270682 243682 270770
rect 243790 270682 243970 270770
rect 244078 270682 244258 270770
rect 244366 270682 244546 270770
rect 244654 270682 244834 270770
rect 244942 270682 245122 270770
rect 245230 270682 245410 270770
rect 245664 270682 245844 270770
rect 245952 270682 246132 270770
rect 246240 270682 246420 270770
rect 246528 270682 246708 270770
rect 246816 270682 246996 270770
rect 247104 270682 247284 270770
rect 247392 270682 247572 270770
rect 247680 270682 247860 270770
rect 248114 270682 248294 270770
rect 248402 270682 248582 270770
rect 248690 270682 248870 270770
rect 248978 270682 249158 270770
rect 249266 270682 249446 270770
rect 249554 270682 249734 270770
rect 249842 270682 250022 270770
rect 250130 270682 250310 270770
rect 250564 270682 250744 270770
rect 360436 270682 360560 270770
rect 360814 270682 360994 270770
rect 361102 270682 361282 270770
rect 361390 270682 361570 270770
rect 361678 270682 361858 270770
rect 361966 270682 362146 270770
rect 362254 270682 362434 270770
rect 362542 270682 362722 270770
rect 362830 270682 363010 270770
rect 363264 270682 363444 270770
rect 363552 270682 363732 270770
rect 363840 270682 364020 270770
rect 364128 270682 364308 270770
rect 364416 270682 364596 270770
rect 364704 270682 364884 270770
rect 364992 270682 365172 270770
rect 365280 270682 365460 270770
rect 365714 270682 365894 270770
rect 366002 270682 366182 270770
rect 366290 270682 366470 270770
rect 366578 270682 366758 270770
rect 366866 270682 367046 270770
rect 367154 270682 367334 270770
rect 367442 270682 367622 270770
rect 367730 270682 367910 270770
rect 243214 270466 243394 270554
rect 243502 270466 243682 270554
rect 243790 270466 243970 270554
rect 244078 270466 244258 270554
rect 244366 270466 244546 270554
rect 244654 270466 244834 270554
rect 244942 270466 245122 270554
rect 245230 270466 245410 270554
rect 245664 270466 245844 270554
rect 245952 270466 246132 270554
rect 246240 270466 246420 270554
rect 246528 270466 246708 270554
rect 246816 270466 246996 270554
rect 247104 270466 247284 270554
rect 247392 270466 247572 270554
rect 247680 270466 247860 270554
rect 248114 270466 248294 270554
rect 248402 270466 248582 270554
rect 248690 270466 248870 270554
rect 248978 270466 249158 270554
rect 249266 270466 249446 270554
rect 249554 270466 249734 270554
rect 249842 270466 250022 270554
rect 250130 270466 250310 270554
rect 250564 270466 250744 270554
rect 360436 270466 360560 270554
rect 360814 270466 360994 270554
rect 361102 270466 361282 270554
rect 361390 270466 361570 270554
rect 361678 270466 361858 270554
rect 361966 270466 362146 270554
rect 362254 270466 362434 270554
rect 362542 270466 362722 270554
rect 362830 270466 363010 270554
rect 363264 270466 363444 270554
rect 363552 270466 363732 270554
rect 363840 270466 364020 270554
rect 364128 270466 364308 270554
rect 364416 270466 364596 270554
rect 364704 270466 364884 270554
rect 364992 270466 365172 270554
rect 365280 270466 365460 270554
rect 365714 270466 365894 270554
rect 366002 270466 366182 270554
rect 366290 270466 366470 270554
rect 366578 270466 366758 270554
rect 366866 270466 367046 270554
rect 367154 270466 367334 270554
rect 367442 270466 367622 270554
rect 367730 270466 367910 270554
rect 243214 269990 243394 270078
rect 243502 269990 243682 270078
rect 243790 269990 243970 270078
rect 244078 269990 244258 270078
rect 244366 269990 244546 270078
rect 244654 269990 244834 270078
rect 244942 269990 245122 270078
rect 245230 269990 245410 270078
rect 245664 269990 245844 270078
rect 245952 269990 246132 270078
rect 246240 269990 246420 270078
rect 246528 269990 246708 270078
rect 246816 269990 246996 270078
rect 247104 269990 247284 270078
rect 247392 269990 247572 270078
rect 247680 269990 247860 270078
rect 248114 269990 248294 270078
rect 248402 269990 248582 270078
rect 248690 269990 248870 270078
rect 248978 269990 249158 270078
rect 249266 269990 249446 270078
rect 249554 269990 249734 270078
rect 249842 269990 250022 270078
rect 250130 269990 250310 270078
rect 250564 269990 250744 270078
rect 360436 269990 360560 270078
rect 360814 269990 360994 270078
rect 361102 269990 361282 270078
rect 361390 269990 361570 270078
rect 361678 269990 361858 270078
rect 361966 269990 362146 270078
rect 362254 269990 362434 270078
rect 362542 269990 362722 270078
rect 362830 269990 363010 270078
rect 363264 269990 363444 270078
rect 363552 269990 363732 270078
rect 363840 269990 364020 270078
rect 364128 269990 364308 270078
rect 364416 269990 364596 270078
rect 364704 269990 364884 270078
rect 364992 269990 365172 270078
rect 365280 269990 365460 270078
rect 365714 269990 365894 270078
rect 366002 269990 366182 270078
rect 366290 269990 366470 270078
rect 366578 269990 366758 270078
rect 366866 269990 367046 270078
rect 367154 269990 367334 270078
rect 367442 269990 367622 270078
rect 367730 269990 367910 270078
rect 243214 269516 243394 269604
rect 243502 269516 243682 269604
rect 243790 269516 243970 269604
rect 244078 269516 244258 269604
rect 244366 269516 244546 269604
rect 244654 269516 244834 269604
rect 244942 269516 245122 269604
rect 245230 269516 245410 269604
rect 245664 269516 245844 269604
rect 245952 269516 246132 269604
rect 246240 269516 246420 269604
rect 246528 269516 246708 269604
rect 246816 269516 246996 269604
rect 247104 269516 247284 269604
rect 247392 269516 247572 269604
rect 247680 269516 247860 269604
rect 248114 269516 248294 269604
rect 248402 269516 248582 269604
rect 248690 269516 248870 269604
rect 248978 269516 249158 269604
rect 249266 269516 249446 269604
rect 249554 269516 249734 269604
rect 249842 269516 250022 269604
rect 250130 269516 250310 269604
rect 250564 269516 250744 269604
rect 360436 269516 360560 269604
rect 360814 269516 360994 269604
rect 361102 269516 361282 269604
rect 361390 269516 361570 269604
rect 361678 269516 361858 269604
rect 361966 269516 362146 269604
rect 362254 269516 362434 269604
rect 362542 269516 362722 269604
rect 362830 269516 363010 269604
rect 363264 269516 363444 269604
rect 363552 269516 363732 269604
rect 363840 269516 364020 269604
rect 364128 269516 364308 269604
rect 364416 269516 364596 269604
rect 364704 269516 364884 269604
rect 364992 269516 365172 269604
rect 365280 269516 365460 269604
rect 365714 269516 365894 269604
rect 366002 269516 366182 269604
rect 366290 269516 366470 269604
rect 366578 269516 366758 269604
rect 366866 269516 367046 269604
rect 367154 269516 367334 269604
rect 367442 269516 367622 269604
rect 367730 269516 367910 269604
rect 243214 269040 243394 269128
rect 243502 269040 243682 269128
rect 243790 269040 243970 269128
rect 244078 269040 244258 269128
rect 244366 269040 244546 269128
rect 244654 269040 244834 269128
rect 244942 269040 245122 269128
rect 245230 269040 245410 269128
rect 245664 269040 245844 269128
rect 245952 269040 246132 269128
rect 246240 269040 246420 269128
rect 246528 269040 246708 269128
rect 246816 269040 246996 269128
rect 247104 269040 247284 269128
rect 247392 269040 247572 269128
rect 247680 269040 247860 269128
rect 248114 269040 248294 269128
rect 248402 269040 248582 269128
rect 248690 269040 248870 269128
rect 248978 269040 249158 269128
rect 249266 269040 249446 269128
rect 249554 269040 249734 269128
rect 249842 269040 250022 269128
rect 250130 269040 250310 269128
rect 250564 269040 250744 269128
rect 360436 269040 360560 269128
rect 360814 269040 360994 269128
rect 361102 269040 361282 269128
rect 361390 269040 361570 269128
rect 361678 269040 361858 269128
rect 361966 269040 362146 269128
rect 362254 269040 362434 269128
rect 362542 269040 362722 269128
rect 362830 269040 363010 269128
rect 363264 269040 363444 269128
rect 363552 269040 363732 269128
rect 363840 269040 364020 269128
rect 364128 269040 364308 269128
rect 364416 269040 364596 269128
rect 364704 269040 364884 269128
rect 364992 269040 365172 269128
rect 365280 269040 365460 269128
rect 365714 269040 365894 269128
rect 366002 269040 366182 269128
rect 366290 269040 366470 269128
rect 366578 269040 366758 269128
rect 366866 269040 367046 269128
rect 367154 269040 367334 269128
rect 367442 269040 367622 269128
rect 367730 269040 367910 269128
rect 243214 268824 243394 268912
rect 243502 268824 243682 268912
rect 243790 268824 243970 268912
rect 244078 268824 244258 268912
rect 244366 268824 244546 268912
rect 244654 268824 244834 268912
rect 244942 268824 245122 268912
rect 245230 268824 245410 268912
rect 245664 268824 245844 268912
rect 245952 268824 246132 268912
rect 246240 268824 246420 268912
rect 246528 268824 246708 268912
rect 246816 268824 246996 268912
rect 247104 268824 247284 268912
rect 247392 268824 247572 268912
rect 247680 268824 247860 268912
rect 248114 268824 248294 268912
rect 248402 268824 248582 268912
rect 248690 268824 248870 268912
rect 248978 268824 249158 268912
rect 249266 268824 249446 268912
rect 249554 268824 249734 268912
rect 249842 268824 250022 268912
rect 250130 268824 250310 268912
rect 250564 268824 250744 268912
rect 360436 268824 360560 268912
rect 360814 268824 360994 268912
rect 361102 268824 361282 268912
rect 361390 268824 361570 268912
rect 361678 268824 361858 268912
rect 361966 268824 362146 268912
rect 362254 268824 362434 268912
rect 362542 268824 362722 268912
rect 362830 268824 363010 268912
rect 363264 268824 363444 268912
rect 363552 268824 363732 268912
rect 363840 268824 364020 268912
rect 364128 268824 364308 268912
rect 364416 268824 364596 268912
rect 364704 268824 364884 268912
rect 364992 268824 365172 268912
rect 365280 268824 365460 268912
rect 365714 268824 365894 268912
rect 366002 268824 366182 268912
rect 366290 268824 366470 268912
rect 366578 268824 366758 268912
rect 366866 268824 367046 268912
rect 367154 268824 367334 268912
rect 367442 268824 367622 268912
rect 367730 268824 367910 268912
rect 243214 268348 243394 268436
rect 243502 268348 243682 268436
rect 243790 268348 243970 268436
rect 244078 268348 244258 268436
rect 244366 268348 244546 268436
rect 244654 268348 244834 268436
rect 244942 268348 245122 268436
rect 245230 268348 245410 268436
rect 245664 268348 245844 268436
rect 245952 268348 246132 268436
rect 246240 268348 246420 268436
rect 246528 268348 246708 268436
rect 246816 268348 246996 268436
rect 247104 268348 247284 268436
rect 247392 268348 247572 268436
rect 247680 268348 247860 268436
rect 248114 268348 248294 268436
rect 248402 268348 248582 268436
rect 248690 268348 248870 268436
rect 248978 268348 249158 268436
rect 249266 268348 249446 268436
rect 249554 268348 249734 268436
rect 249842 268348 250022 268436
rect 250130 268348 250310 268436
rect 250564 268348 250744 268436
rect 360436 268348 360560 268436
rect 360814 268348 360994 268436
rect 361102 268348 361282 268436
rect 361390 268348 361570 268436
rect 361678 268348 361858 268436
rect 361966 268348 362146 268436
rect 362254 268348 362434 268436
rect 362542 268348 362722 268436
rect 362830 268348 363010 268436
rect 363264 268348 363444 268436
rect 363552 268348 363732 268436
rect 363840 268348 364020 268436
rect 364128 268348 364308 268436
rect 364416 268348 364596 268436
rect 364704 268348 364884 268436
rect 364992 268348 365172 268436
rect 365280 268348 365460 268436
rect 365714 268348 365894 268436
rect 366002 268348 366182 268436
rect 366290 268348 366470 268436
rect 366578 268348 366758 268436
rect 366866 268348 367046 268436
rect 367154 268348 367334 268436
rect 367442 268348 367622 268436
rect 367730 268348 367910 268436
rect 243214 268132 243394 268220
rect 243502 268132 243682 268220
rect 243790 268132 243970 268220
rect 244078 268132 244258 268220
rect 244366 268132 244546 268220
rect 244654 268132 244834 268220
rect 244942 268132 245122 268220
rect 245230 268132 245410 268220
rect 245664 268132 245844 268220
rect 245952 268132 246132 268220
rect 246240 268132 246420 268220
rect 246528 268132 246708 268220
rect 246816 268132 246996 268220
rect 247104 268132 247284 268220
rect 247392 268132 247572 268220
rect 247680 268132 247860 268220
rect 248114 268132 248294 268220
rect 248402 268132 248582 268220
rect 248690 268132 248870 268220
rect 248978 268132 249158 268220
rect 249266 268132 249446 268220
rect 249554 268132 249734 268220
rect 249842 268132 250022 268220
rect 250130 268132 250310 268220
rect 250564 268132 250744 268220
rect 360436 268132 360560 268220
rect 360814 268132 360994 268220
rect 361102 268132 361282 268220
rect 361390 268132 361570 268220
rect 361678 268132 361858 268220
rect 361966 268132 362146 268220
rect 362254 268132 362434 268220
rect 362542 268132 362722 268220
rect 362830 268132 363010 268220
rect 363264 268132 363444 268220
rect 363552 268132 363732 268220
rect 363840 268132 364020 268220
rect 364128 268132 364308 268220
rect 364416 268132 364596 268220
rect 364704 268132 364884 268220
rect 364992 268132 365172 268220
rect 365280 268132 365460 268220
rect 365714 268132 365894 268220
rect 366002 268132 366182 268220
rect 366290 268132 366470 268220
rect 366578 268132 366758 268220
rect 366866 268132 367046 268220
rect 367154 268132 367334 268220
rect 367442 268132 367622 268220
rect 367730 268132 367910 268220
rect 243214 267656 243394 267744
rect 243502 267656 243682 267744
rect 243790 267656 243970 267744
rect 244078 267656 244258 267744
rect 244366 267656 244546 267744
rect 244654 267656 244834 267744
rect 244942 267656 245122 267744
rect 245230 267656 245410 267744
rect 245664 267656 245844 267744
rect 245952 267656 246132 267744
rect 246240 267656 246420 267744
rect 246528 267656 246708 267744
rect 246816 267656 246996 267744
rect 247104 267656 247284 267744
rect 247392 267656 247572 267744
rect 247680 267656 247860 267744
rect 248114 267656 248294 267744
rect 248402 267656 248582 267744
rect 248690 267656 248870 267744
rect 248978 267656 249158 267744
rect 249266 267656 249446 267744
rect 249554 267656 249734 267744
rect 249842 267656 250022 267744
rect 250130 267656 250310 267744
rect 250564 267656 250744 267744
rect 360436 267656 360560 267744
rect 360814 267656 360994 267744
rect 361102 267656 361282 267744
rect 361390 267656 361570 267744
rect 361678 267656 361858 267744
rect 361966 267656 362146 267744
rect 362254 267656 362434 267744
rect 362542 267656 362722 267744
rect 362830 267656 363010 267744
rect 363264 267656 363444 267744
rect 363552 267656 363732 267744
rect 363840 267656 364020 267744
rect 364128 267656 364308 267744
rect 364416 267656 364596 267744
rect 364704 267656 364884 267744
rect 364992 267656 365172 267744
rect 365280 267656 365460 267744
rect 365714 267656 365894 267744
rect 366002 267656 366182 267744
rect 366290 267656 366470 267744
rect 366578 267656 366758 267744
rect 366866 267656 367046 267744
rect 367154 267656 367334 267744
rect 367442 267656 367622 267744
rect 367730 267656 367910 267744
rect 243214 267440 243394 267528
rect 243502 267440 243682 267528
rect 243790 267440 243970 267528
rect 244078 267440 244258 267528
rect 244366 267440 244546 267528
rect 244654 267440 244834 267528
rect 244942 267440 245122 267528
rect 245230 267440 245410 267528
rect 245664 267440 245844 267528
rect 245952 267440 246132 267528
rect 246240 267440 246420 267528
rect 246528 267440 246708 267528
rect 246816 267440 246996 267528
rect 247104 267440 247284 267528
rect 247392 267440 247572 267528
rect 247680 267440 247860 267528
rect 248114 267440 248294 267528
rect 248402 267440 248582 267528
rect 248690 267440 248870 267528
rect 248978 267440 249158 267528
rect 249266 267440 249446 267528
rect 249554 267440 249734 267528
rect 249842 267440 250022 267528
rect 250130 267440 250310 267528
rect 250564 267440 250744 267528
rect 360436 267440 360560 267528
rect 360814 267440 360994 267528
rect 361102 267440 361282 267528
rect 361390 267440 361570 267528
rect 361678 267440 361858 267528
rect 361966 267440 362146 267528
rect 362254 267440 362434 267528
rect 362542 267440 362722 267528
rect 362830 267440 363010 267528
rect 363264 267440 363444 267528
rect 363552 267440 363732 267528
rect 363840 267440 364020 267528
rect 364128 267440 364308 267528
rect 364416 267440 364596 267528
rect 364704 267440 364884 267528
rect 364992 267440 365172 267528
rect 365280 267440 365460 267528
rect 365714 267440 365894 267528
rect 366002 267440 366182 267528
rect 366290 267440 366470 267528
rect 366578 267440 366758 267528
rect 366866 267440 367046 267528
rect 367154 267440 367334 267528
rect 367442 267440 367622 267528
rect 367730 267440 367910 267528
rect 243214 266964 243394 267052
rect 243502 266964 243682 267052
rect 243790 266964 243970 267052
rect 244078 266964 244258 267052
rect 244366 266964 244546 267052
rect 244654 266964 244834 267052
rect 244942 266964 245122 267052
rect 245230 266964 245410 267052
rect 245664 266964 245844 267052
rect 245952 266964 246132 267052
rect 246240 266964 246420 267052
rect 246528 266964 246708 267052
rect 246816 266964 246996 267052
rect 247104 266964 247284 267052
rect 247392 266964 247572 267052
rect 247680 266964 247860 267052
rect 248114 266964 248294 267052
rect 248402 266964 248582 267052
rect 248690 266964 248870 267052
rect 248978 266964 249158 267052
rect 249266 266964 249446 267052
rect 249554 266964 249734 267052
rect 249842 266964 250022 267052
rect 250130 266964 250310 267052
rect 250564 266964 250744 267052
rect 360436 266964 360560 267052
rect 360814 266964 360994 267052
rect 361102 266964 361282 267052
rect 361390 266964 361570 267052
rect 361678 266964 361858 267052
rect 361966 266964 362146 267052
rect 362254 266964 362434 267052
rect 362542 266964 362722 267052
rect 362830 266964 363010 267052
rect 363264 266964 363444 267052
rect 363552 266964 363732 267052
rect 363840 266964 364020 267052
rect 364128 266964 364308 267052
rect 364416 266964 364596 267052
rect 364704 266964 364884 267052
rect 364992 266964 365172 267052
rect 365280 266964 365460 267052
rect 365714 266964 365894 267052
rect 366002 266964 366182 267052
rect 366290 266964 366470 267052
rect 366578 266964 366758 267052
rect 366866 266964 367046 267052
rect 367154 266964 367334 267052
rect 367442 266964 367622 267052
rect 367730 266964 367910 267052
rect 243214 266490 243394 266578
rect 243502 266490 243682 266578
rect 243790 266490 243970 266578
rect 244078 266490 244258 266578
rect 244366 266490 244546 266578
rect 244654 266490 244834 266578
rect 244942 266490 245122 266578
rect 245230 266490 245410 266578
rect 245664 266490 245844 266578
rect 245952 266490 246132 266578
rect 246240 266490 246420 266578
rect 246528 266490 246708 266578
rect 246816 266490 246996 266578
rect 247104 266490 247284 266578
rect 247392 266490 247572 266578
rect 247680 266490 247860 266578
rect 248114 266490 248294 266578
rect 248402 266490 248582 266578
rect 248690 266490 248870 266578
rect 248978 266490 249158 266578
rect 249266 266490 249446 266578
rect 249554 266490 249734 266578
rect 249842 266490 250022 266578
rect 250130 266490 250310 266578
rect 250564 266490 250744 266578
rect 360436 266490 360560 266578
rect 360814 266490 360994 266578
rect 361102 266490 361282 266578
rect 361390 266490 361570 266578
rect 361678 266490 361858 266578
rect 361966 266490 362146 266578
rect 362254 266490 362434 266578
rect 362542 266490 362722 266578
rect 362830 266490 363010 266578
rect 363264 266490 363444 266578
rect 363552 266490 363732 266578
rect 363840 266490 364020 266578
rect 364128 266490 364308 266578
rect 364416 266490 364596 266578
rect 364704 266490 364884 266578
rect 364992 266490 365172 266578
rect 365280 266490 365460 266578
rect 365714 266490 365894 266578
rect 366002 266490 366182 266578
rect 366290 266490 366470 266578
rect 366578 266490 366758 266578
rect 366866 266490 367046 266578
rect 367154 266490 367334 266578
rect 367442 266490 367622 266578
rect 367730 266490 367910 266578
rect 243214 266014 243394 266102
rect 243502 266014 243682 266102
rect 243790 266014 243970 266102
rect 244078 266014 244258 266102
rect 244366 266014 244546 266102
rect 244654 266014 244834 266102
rect 244942 266014 245122 266102
rect 245230 266014 245410 266102
rect 245664 266014 245844 266102
rect 245952 266014 246132 266102
rect 246240 266014 246420 266102
rect 246528 266014 246708 266102
rect 246816 266014 246996 266102
rect 247104 266014 247284 266102
rect 247392 266014 247572 266102
rect 247680 266014 247860 266102
rect 248114 266014 248294 266102
rect 248402 266014 248582 266102
rect 248690 266014 248870 266102
rect 248978 266014 249158 266102
rect 249266 266014 249446 266102
rect 249554 266014 249734 266102
rect 249842 266014 250022 266102
rect 250130 266014 250310 266102
rect 250564 266014 250744 266102
rect 360436 266014 360560 266102
rect 360814 266014 360994 266102
rect 361102 266014 361282 266102
rect 361390 266014 361570 266102
rect 361678 266014 361858 266102
rect 361966 266014 362146 266102
rect 362254 266014 362434 266102
rect 362542 266014 362722 266102
rect 362830 266014 363010 266102
rect 363264 266014 363444 266102
rect 363552 266014 363732 266102
rect 363840 266014 364020 266102
rect 364128 266014 364308 266102
rect 364416 266014 364596 266102
rect 364704 266014 364884 266102
rect 364992 266014 365172 266102
rect 365280 266014 365460 266102
rect 365714 266014 365894 266102
rect 366002 266014 366182 266102
rect 366290 266014 366470 266102
rect 366578 266014 366758 266102
rect 366866 266014 367046 266102
rect 367154 266014 367334 266102
rect 367442 266014 367622 266102
rect 367730 266014 367910 266102
rect 243214 265798 243394 265886
rect 243502 265798 243682 265886
rect 243790 265798 243970 265886
rect 244078 265798 244258 265886
rect 244366 265798 244546 265886
rect 244654 265798 244834 265886
rect 244942 265798 245122 265886
rect 245230 265798 245410 265886
rect 245664 265798 245844 265886
rect 245952 265798 246132 265886
rect 246240 265798 246420 265886
rect 246528 265798 246708 265886
rect 246816 265798 246996 265886
rect 247104 265798 247284 265886
rect 247392 265798 247572 265886
rect 247680 265798 247860 265886
rect 248114 265798 248294 265886
rect 248402 265798 248582 265886
rect 248690 265798 248870 265886
rect 248978 265798 249158 265886
rect 249266 265798 249446 265886
rect 249554 265798 249734 265886
rect 249842 265798 250022 265886
rect 250130 265798 250310 265886
rect 250564 265798 250744 265886
rect 360436 265798 360560 265886
rect 360814 265798 360994 265886
rect 361102 265798 361282 265886
rect 361390 265798 361570 265886
rect 361678 265798 361858 265886
rect 361966 265798 362146 265886
rect 362254 265798 362434 265886
rect 362542 265798 362722 265886
rect 362830 265798 363010 265886
rect 363264 265798 363444 265886
rect 363552 265798 363732 265886
rect 363840 265798 364020 265886
rect 364128 265798 364308 265886
rect 364416 265798 364596 265886
rect 364704 265798 364884 265886
rect 364992 265798 365172 265886
rect 365280 265798 365460 265886
rect 365714 265798 365894 265886
rect 366002 265798 366182 265886
rect 366290 265798 366470 265886
rect 366578 265798 366758 265886
rect 366866 265798 367046 265886
rect 367154 265798 367334 265886
rect 367442 265798 367622 265886
rect 367730 265798 367910 265886
rect 243214 265322 243394 265410
rect 243502 265322 243682 265410
rect 243790 265322 243970 265410
rect 244078 265322 244258 265410
rect 244366 265322 244546 265410
rect 244654 265322 244834 265410
rect 244942 265322 245122 265410
rect 245230 265322 245410 265410
rect 245664 265322 245844 265410
rect 245952 265322 246132 265410
rect 246240 265322 246420 265410
rect 246528 265322 246708 265410
rect 246816 265322 246996 265410
rect 247104 265322 247284 265410
rect 247392 265322 247572 265410
rect 247680 265322 247860 265410
rect 248114 265322 248294 265410
rect 248402 265322 248582 265410
rect 248690 265322 248870 265410
rect 248978 265322 249158 265410
rect 249266 265322 249446 265410
rect 249554 265322 249734 265410
rect 249842 265322 250022 265410
rect 250130 265322 250310 265410
rect 250564 265322 250744 265410
rect 360436 265322 360560 265410
rect 360814 265322 360994 265410
rect 361102 265322 361282 265410
rect 361390 265322 361570 265410
rect 361678 265322 361858 265410
rect 361966 265322 362146 265410
rect 362254 265322 362434 265410
rect 362542 265322 362722 265410
rect 362830 265322 363010 265410
rect 363264 265322 363444 265410
rect 363552 265322 363732 265410
rect 363840 265322 364020 265410
rect 364128 265322 364308 265410
rect 364416 265322 364596 265410
rect 364704 265322 364884 265410
rect 364992 265322 365172 265410
rect 365280 265322 365460 265410
rect 365714 265322 365894 265410
rect 366002 265322 366182 265410
rect 366290 265322 366470 265410
rect 366578 265322 366758 265410
rect 366866 265322 367046 265410
rect 367154 265322 367334 265410
rect 367442 265322 367622 265410
rect 367730 265322 367910 265410
rect 243214 265106 243394 265194
rect 243502 265106 243682 265194
rect 243790 265106 243970 265194
rect 244078 265106 244258 265194
rect 244366 265106 244546 265194
rect 244654 265106 244834 265194
rect 244942 265106 245122 265194
rect 245230 265106 245410 265194
rect 245664 265106 245844 265194
rect 245952 265106 246132 265194
rect 246240 265106 246420 265194
rect 246528 265106 246708 265194
rect 246816 265106 246996 265194
rect 247104 265106 247284 265194
rect 247392 265106 247572 265194
rect 247680 265106 247860 265194
rect 248114 265106 248294 265194
rect 248402 265106 248582 265194
rect 248690 265106 248870 265194
rect 248978 265106 249158 265194
rect 249266 265106 249446 265194
rect 249554 265106 249734 265194
rect 249842 265106 250022 265194
rect 250130 265106 250310 265194
rect 250564 265106 250744 265194
rect 360436 265106 360560 265194
rect 360814 265106 360994 265194
rect 361102 265106 361282 265194
rect 361390 265106 361570 265194
rect 361678 265106 361858 265194
rect 361966 265106 362146 265194
rect 362254 265106 362434 265194
rect 362542 265106 362722 265194
rect 362830 265106 363010 265194
rect 363264 265106 363444 265194
rect 363552 265106 363732 265194
rect 363840 265106 364020 265194
rect 364128 265106 364308 265194
rect 364416 265106 364596 265194
rect 364704 265106 364884 265194
rect 364992 265106 365172 265194
rect 365280 265106 365460 265194
rect 365714 265106 365894 265194
rect 366002 265106 366182 265194
rect 366290 265106 366470 265194
rect 366578 265106 366758 265194
rect 366866 265106 367046 265194
rect 367154 265106 367334 265194
rect 367442 265106 367622 265194
rect 367730 265106 367910 265194
rect 243214 264630 243394 264718
rect 243502 264630 243682 264718
rect 243790 264630 243970 264718
rect 244078 264630 244258 264718
rect 244366 264630 244546 264718
rect 244654 264630 244834 264718
rect 244942 264630 245122 264718
rect 245230 264630 245410 264718
rect 245664 264630 245844 264718
rect 245952 264630 246132 264718
rect 246240 264630 246420 264718
rect 246528 264630 246708 264718
rect 246816 264630 246996 264718
rect 247104 264630 247284 264718
rect 247392 264630 247572 264718
rect 247680 264630 247860 264718
rect 248114 264630 248294 264718
rect 248402 264630 248582 264718
rect 248690 264630 248870 264718
rect 248978 264630 249158 264718
rect 249266 264630 249446 264718
rect 249554 264630 249734 264718
rect 249842 264630 250022 264718
rect 250130 264630 250310 264718
rect 250564 264630 250744 264718
rect 360436 264630 360560 264718
rect 360814 264630 360994 264718
rect 361102 264630 361282 264718
rect 361390 264630 361570 264718
rect 361678 264630 361858 264718
rect 361966 264630 362146 264718
rect 362254 264630 362434 264718
rect 362542 264630 362722 264718
rect 362830 264630 363010 264718
rect 363264 264630 363444 264718
rect 363552 264630 363732 264718
rect 363840 264630 364020 264718
rect 364128 264630 364308 264718
rect 364416 264630 364596 264718
rect 364704 264630 364884 264718
rect 364992 264630 365172 264718
rect 365280 264630 365460 264718
rect 365714 264630 365894 264718
rect 366002 264630 366182 264718
rect 366290 264630 366470 264718
rect 366578 264630 366758 264718
rect 366866 264630 367046 264718
rect 367154 264630 367334 264718
rect 367442 264630 367622 264718
rect 367730 264630 367910 264718
rect 243214 264414 243394 264502
rect 243502 264414 243682 264502
rect 243790 264414 243970 264502
rect 244078 264414 244258 264502
rect 244366 264414 244546 264502
rect 244654 264414 244834 264502
rect 244942 264414 245122 264502
rect 245230 264414 245410 264502
rect 245664 264414 245844 264502
rect 245952 264414 246132 264502
rect 246240 264414 246420 264502
rect 246528 264414 246708 264502
rect 246816 264414 246996 264502
rect 247104 264414 247284 264502
rect 247392 264414 247572 264502
rect 247680 264414 247860 264502
rect 248114 264414 248294 264502
rect 248402 264414 248582 264502
rect 248690 264414 248870 264502
rect 248978 264414 249158 264502
rect 249266 264414 249446 264502
rect 249554 264414 249734 264502
rect 249842 264414 250022 264502
rect 250130 264414 250310 264502
rect 250564 264414 250744 264502
rect 360436 264414 360560 264502
rect 360814 264414 360994 264502
rect 361102 264414 361282 264502
rect 361390 264414 361570 264502
rect 361678 264414 361858 264502
rect 361966 264414 362146 264502
rect 362254 264414 362434 264502
rect 362542 264414 362722 264502
rect 362830 264414 363010 264502
rect 363264 264414 363444 264502
rect 363552 264414 363732 264502
rect 363840 264414 364020 264502
rect 364128 264414 364308 264502
rect 364416 264414 364596 264502
rect 364704 264414 364884 264502
rect 364992 264414 365172 264502
rect 365280 264414 365460 264502
rect 365714 264414 365894 264502
rect 366002 264414 366182 264502
rect 366290 264414 366470 264502
rect 366578 264414 366758 264502
rect 366866 264414 367046 264502
rect 367154 264414 367334 264502
rect 367442 264414 367622 264502
rect 367730 264414 367910 264502
rect 243214 263938 243394 264026
rect 243502 263938 243682 264026
rect 243790 263938 243970 264026
rect 244078 263938 244258 264026
rect 244366 263938 244546 264026
rect 244654 263938 244834 264026
rect 244942 263938 245122 264026
rect 245230 263938 245410 264026
rect 245664 263938 245844 264026
rect 245952 263938 246132 264026
rect 246240 263938 246420 264026
rect 246528 263938 246708 264026
rect 246816 263938 246996 264026
rect 247104 263938 247284 264026
rect 247392 263938 247572 264026
rect 247680 263938 247860 264026
rect 248114 263938 248294 264026
rect 248402 263938 248582 264026
rect 248690 263938 248870 264026
rect 248978 263938 249158 264026
rect 249266 263938 249446 264026
rect 249554 263938 249734 264026
rect 249842 263938 250022 264026
rect 250130 263938 250310 264026
rect 250564 263938 250744 264026
rect 360436 263938 360560 264026
rect 360814 263938 360994 264026
rect 361102 263938 361282 264026
rect 361390 263938 361570 264026
rect 361678 263938 361858 264026
rect 361966 263938 362146 264026
rect 362254 263938 362434 264026
rect 362542 263938 362722 264026
rect 362830 263938 363010 264026
rect 363264 263938 363444 264026
rect 363552 263938 363732 264026
rect 363840 263938 364020 264026
rect 364128 263938 364308 264026
rect 364416 263938 364596 264026
rect 364704 263938 364884 264026
rect 364992 263938 365172 264026
rect 365280 263938 365460 264026
rect 365714 263938 365894 264026
rect 366002 263938 366182 264026
rect 366290 263938 366470 264026
rect 366578 263938 366758 264026
rect 366866 263938 367046 264026
rect 367154 263938 367334 264026
rect 367442 263938 367622 264026
rect 367730 263938 367910 264026
rect 243214 263464 243394 263552
rect 243502 263464 243682 263552
rect 243790 263464 243970 263552
rect 244078 263464 244258 263552
rect 244366 263464 244546 263552
rect 244654 263464 244834 263552
rect 244942 263464 245122 263552
rect 245230 263464 245410 263552
rect 245664 263464 245844 263552
rect 245952 263464 246132 263552
rect 246240 263464 246420 263552
rect 246528 263464 246708 263552
rect 246816 263464 246996 263552
rect 247104 263464 247284 263552
rect 247392 263464 247572 263552
rect 247680 263464 247860 263552
rect 248114 263464 248294 263552
rect 248402 263464 248582 263552
rect 248690 263464 248870 263552
rect 248978 263464 249158 263552
rect 249266 263464 249446 263552
rect 249554 263464 249734 263552
rect 249842 263464 250022 263552
rect 250130 263464 250310 263552
rect 250564 263464 250744 263552
rect 360436 263464 360560 263552
rect 360814 263464 360994 263552
rect 361102 263464 361282 263552
rect 361390 263464 361570 263552
rect 361678 263464 361858 263552
rect 361966 263464 362146 263552
rect 362254 263464 362434 263552
rect 362542 263464 362722 263552
rect 362830 263464 363010 263552
rect 363264 263464 363444 263552
rect 363552 263464 363732 263552
rect 363840 263464 364020 263552
rect 364128 263464 364308 263552
rect 364416 263464 364596 263552
rect 364704 263464 364884 263552
rect 364992 263464 365172 263552
rect 365280 263464 365460 263552
rect 365714 263464 365894 263552
rect 366002 263464 366182 263552
rect 366290 263464 366470 263552
rect 366578 263464 366758 263552
rect 366866 263464 367046 263552
rect 367154 263464 367334 263552
rect 367442 263464 367622 263552
rect 367730 263464 367910 263552
rect 243214 262988 243394 263076
rect 243502 262988 243682 263076
rect 243790 262988 243970 263076
rect 244078 262988 244258 263076
rect 244366 262988 244546 263076
rect 244654 262988 244834 263076
rect 244942 262988 245122 263076
rect 245230 262988 245410 263076
rect 245664 262988 245844 263076
rect 245952 262988 246132 263076
rect 246240 262988 246420 263076
rect 246528 262988 246708 263076
rect 246816 262988 246996 263076
rect 247104 262988 247284 263076
rect 247392 262988 247572 263076
rect 247680 262988 247860 263076
rect 248114 262988 248294 263076
rect 248402 262988 248582 263076
rect 248690 262988 248870 263076
rect 248978 262988 249158 263076
rect 249266 262988 249446 263076
rect 249554 262988 249734 263076
rect 249842 262988 250022 263076
rect 250130 262988 250310 263076
rect 250564 262988 250744 263076
rect 360436 262988 360560 263076
rect 360814 262988 360994 263076
rect 361102 262988 361282 263076
rect 361390 262988 361570 263076
rect 361678 262988 361858 263076
rect 361966 262988 362146 263076
rect 362254 262988 362434 263076
rect 362542 262988 362722 263076
rect 362830 262988 363010 263076
rect 363264 262988 363444 263076
rect 363552 262988 363732 263076
rect 363840 262988 364020 263076
rect 364128 262988 364308 263076
rect 364416 262988 364596 263076
rect 364704 262988 364884 263076
rect 364992 262988 365172 263076
rect 365280 262988 365460 263076
rect 365714 262988 365894 263076
rect 366002 262988 366182 263076
rect 366290 262988 366470 263076
rect 366578 262988 366758 263076
rect 366866 262988 367046 263076
rect 367154 262988 367334 263076
rect 367442 262988 367622 263076
rect 367730 262988 367910 263076
rect 243214 262772 243394 262860
rect 243502 262772 243682 262860
rect 243790 262772 243970 262860
rect 244078 262772 244258 262860
rect 244366 262772 244546 262860
rect 244654 262772 244834 262860
rect 244942 262772 245122 262860
rect 245230 262772 245410 262860
rect 245664 262772 245844 262860
rect 245952 262772 246132 262860
rect 246240 262772 246420 262860
rect 246528 262772 246708 262860
rect 246816 262772 246996 262860
rect 247104 262772 247284 262860
rect 247392 262772 247572 262860
rect 247680 262772 247860 262860
rect 248114 262772 248294 262860
rect 248402 262772 248582 262860
rect 248690 262772 248870 262860
rect 248978 262772 249158 262860
rect 249266 262772 249446 262860
rect 249554 262772 249734 262860
rect 249842 262772 250022 262860
rect 250130 262772 250310 262860
rect 250564 262772 250744 262860
rect 360436 262772 360560 262860
rect 360814 262772 360994 262860
rect 361102 262772 361282 262860
rect 361390 262772 361570 262860
rect 361678 262772 361858 262860
rect 361966 262772 362146 262860
rect 362254 262772 362434 262860
rect 362542 262772 362722 262860
rect 362830 262772 363010 262860
rect 363264 262772 363444 262860
rect 363552 262772 363732 262860
rect 363840 262772 364020 262860
rect 364128 262772 364308 262860
rect 364416 262772 364596 262860
rect 364704 262772 364884 262860
rect 364992 262772 365172 262860
rect 365280 262772 365460 262860
rect 365714 262772 365894 262860
rect 366002 262772 366182 262860
rect 366290 262772 366470 262860
rect 366578 262772 366758 262860
rect 366866 262772 367046 262860
rect 367154 262772 367334 262860
rect 367442 262772 367622 262860
rect 367730 262772 367910 262860
rect 243214 262296 243394 262384
rect 243502 262296 243682 262384
rect 243790 262296 243970 262384
rect 244078 262296 244258 262384
rect 244366 262296 244546 262384
rect 244654 262296 244834 262384
rect 244942 262296 245122 262384
rect 245230 262296 245410 262384
rect 245664 262296 245844 262384
rect 245952 262296 246132 262384
rect 246240 262296 246420 262384
rect 246528 262296 246708 262384
rect 246816 262296 246996 262384
rect 247104 262296 247284 262384
rect 247392 262296 247572 262384
rect 247680 262296 247860 262384
rect 248114 262296 248294 262384
rect 248402 262296 248582 262384
rect 248690 262296 248870 262384
rect 248978 262296 249158 262384
rect 249266 262296 249446 262384
rect 249554 262296 249734 262384
rect 249842 262296 250022 262384
rect 250130 262296 250310 262384
rect 250564 262296 250744 262384
rect 360436 262296 360560 262384
rect 360814 262296 360994 262384
rect 361102 262296 361282 262384
rect 361390 262296 361570 262384
rect 361678 262296 361858 262384
rect 361966 262296 362146 262384
rect 362254 262296 362434 262384
rect 362542 262296 362722 262384
rect 362830 262296 363010 262384
rect 363264 262296 363444 262384
rect 363552 262296 363732 262384
rect 363840 262296 364020 262384
rect 364128 262296 364308 262384
rect 364416 262296 364596 262384
rect 364704 262296 364884 262384
rect 364992 262296 365172 262384
rect 365280 262296 365460 262384
rect 365714 262296 365894 262384
rect 366002 262296 366182 262384
rect 366290 262296 366470 262384
rect 366578 262296 366758 262384
rect 366866 262296 367046 262384
rect 367154 262296 367334 262384
rect 367442 262296 367622 262384
rect 367730 262296 367910 262384
rect 243214 262080 243394 262168
rect 243502 262080 243682 262168
rect 243790 262080 243970 262168
rect 244078 262080 244258 262168
rect 244366 262080 244546 262168
rect 244654 262080 244834 262168
rect 244942 262080 245122 262168
rect 245230 262080 245410 262168
rect 245664 262080 245844 262168
rect 245952 262080 246132 262168
rect 246240 262080 246420 262168
rect 246528 262080 246708 262168
rect 246816 262080 246996 262168
rect 247104 262080 247284 262168
rect 247392 262080 247572 262168
rect 247680 262080 247860 262168
rect 248114 262080 248294 262168
rect 248402 262080 248582 262168
rect 248690 262080 248870 262168
rect 248978 262080 249158 262168
rect 249266 262080 249446 262168
rect 249554 262080 249734 262168
rect 249842 262080 250022 262168
rect 250130 262080 250310 262168
rect 250564 262080 250744 262168
rect 360436 262080 360560 262168
rect 360814 262080 360994 262168
rect 361102 262080 361282 262168
rect 361390 262080 361570 262168
rect 361678 262080 361858 262168
rect 361966 262080 362146 262168
rect 362254 262080 362434 262168
rect 362542 262080 362722 262168
rect 362830 262080 363010 262168
rect 363264 262080 363444 262168
rect 363552 262080 363732 262168
rect 363840 262080 364020 262168
rect 364128 262080 364308 262168
rect 364416 262080 364596 262168
rect 364704 262080 364884 262168
rect 364992 262080 365172 262168
rect 365280 262080 365460 262168
rect 365714 262080 365894 262168
rect 366002 262080 366182 262168
rect 366290 262080 366470 262168
rect 366578 262080 366758 262168
rect 366866 262080 367046 262168
rect 367154 262080 367334 262168
rect 367442 262080 367622 262168
rect 367730 262080 367910 262168
rect 243214 261604 243394 261692
rect 243502 261604 243682 261692
rect 243790 261604 243970 261692
rect 244078 261604 244258 261692
rect 244366 261604 244546 261692
rect 244654 261604 244834 261692
rect 244942 261604 245122 261692
rect 245230 261604 245410 261692
rect 245664 261604 245844 261692
rect 245952 261604 246132 261692
rect 246240 261604 246420 261692
rect 246528 261604 246708 261692
rect 246816 261604 246996 261692
rect 247104 261604 247284 261692
rect 247392 261604 247572 261692
rect 247680 261604 247860 261692
rect 248114 261604 248294 261692
rect 248402 261604 248582 261692
rect 248690 261604 248870 261692
rect 248978 261604 249158 261692
rect 249266 261604 249446 261692
rect 249554 261604 249734 261692
rect 249842 261604 250022 261692
rect 250130 261604 250310 261692
rect 250564 261604 250744 261692
rect 360436 261604 360560 261692
rect 360814 261604 360994 261692
rect 361102 261604 361282 261692
rect 361390 261604 361570 261692
rect 361678 261604 361858 261692
rect 361966 261604 362146 261692
rect 362254 261604 362434 261692
rect 362542 261604 362722 261692
rect 362830 261604 363010 261692
rect 363264 261604 363444 261692
rect 363552 261604 363732 261692
rect 363840 261604 364020 261692
rect 364128 261604 364308 261692
rect 364416 261604 364596 261692
rect 364704 261604 364884 261692
rect 364992 261604 365172 261692
rect 365280 261604 365460 261692
rect 365714 261604 365894 261692
rect 366002 261604 366182 261692
rect 366290 261604 366470 261692
rect 366578 261604 366758 261692
rect 366866 261604 367046 261692
rect 367154 261604 367334 261692
rect 367442 261604 367622 261692
rect 367730 261604 367910 261692
rect 243214 261388 243394 261476
rect 243502 261388 243682 261476
rect 243790 261388 243970 261476
rect 244078 261388 244258 261476
rect 244366 261388 244546 261476
rect 244654 261388 244834 261476
rect 244942 261388 245122 261476
rect 245230 261388 245410 261476
rect 245664 261388 245844 261476
rect 245952 261388 246132 261476
rect 246240 261388 246420 261476
rect 246528 261388 246708 261476
rect 246816 261388 246996 261476
rect 247104 261388 247284 261476
rect 247392 261388 247572 261476
rect 247680 261388 247860 261476
rect 248114 261388 248294 261476
rect 248402 261388 248582 261476
rect 248690 261388 248870 261476
rect 248978 261388 249158 261476
rect 249266 261388 249446 261476
rect 249554 261388 249734 261476
rect 249842 261388 250022 261476
rect 250130 261388 250310 261476
rect 250564 261388 250744 261476
rect 360436 261388 360560 261476
rect 360814 261388 360994 261476
rect 361102 261388 361282 261476
rect 361390 261388 361570 261476
rect 361678 261388 361858 261476
rect 361966 261388 362146 261476
rect 362254 261388 362434 261476
rect 362542 261388 362722 261476
rect 362830 261388 363010 261476
rect 363264 261388 363444 261476
rect 363552 261388 363732 261476
rect 363840 261388 364020 261476
rect 364128 261388 364308 261476
rect 364416 261388 364596 261476
rect 364704 261388 364884 261476
rect 364992 261388 365172 261476
rect 365280 261388 365460 261476
rect 365714 261388 365894 261476
rect 366002 261388 366182 261476
rect 366290 261388 366470 261476
rect 366578 261388 366758 261476
rect 366866 261388 367046 261476
rect 367154 261388 367334 261476
rect 367442 261388 367622 261476
rect 367730 261388 367910 261476
rect 243214 260912 243394 261000
rect 243502 260912 243682 261000
rect 243790 260912 243970 261000
rect 244078 260912 244258 261000
rect 244366 260912 244546 261000
rect 244654 260912 244834 261000
rect 244942 260912 245122 261000
rect 245230 260912 245410 261000
rect 245664 260912 245844 261000
rect 245952 260912 246132 261000
rect 246240 260912 246420 261000
rect 246528 260912 246708 261000
rect 246816 260912 246996 261000
rect 247104 260912 247284 261000
rect 247392 260912 247572 261000
rect 247680 260912 247860 261000
rect 248114 260912 248294 261000
rect 248402 260912 248582 261000
rect 248690 260912 248870 261000
rect 248978 260912 249158 261000
rect 249266 260912 249446 261000
rect 249554 260912 249734 261000
rect 249842 260912 250022 261000
rect 250130 260912 250310 261000
rect 250564 260912 250744 261000
rect 360436 260912 360560 261000
rect 360814 260912 360994 261000
rect 361102 260912 361282 261000
rect 361390 260912 361570 261000
rect 361678 260912 361858 261000
rect 361966 260912 362146 261000
rect 362254 260912 362434 261000
rect 362542 260912 362722 261000
rect 362830 260912 363010 261000
rect 363264 260912 363444 261000
rect 363552 260912 363732 261000
rect 363840 260912 364020 261000
rect 364128 260912 364308 261000
rect 364416 260912 364596 261000
rect 364704 260912 364884 261000
rect 364992 260912 365172 261000
rect 365280 260912 365460 261000
rect 365714 260912 365894 261000
rect 366002 260912 366182 261000
rect 366290 260912 366470 261000
rect 366578 260912 366758 261000
rect 366866 260912 367046 261000
rect 367154 260912 367334 261000
rect 367442 260912 367622 261000
rect 367730 260912 367910 261000
rect 243214 260438 243394 260526
rect 243502 260438 243682 260526
rect 243790 260438 243970 260526
rect 244078 260438 244258 260526
rect 244366 260438 244546 260526
rect 244654 260438 244834 260526
rect 244942 260438 245122 260526
rect 245230 260438 245410 260526
rect 245664 260438 245844 260526
rect 245952 260438 246132 260526
rect 246240 260438 246420 260526
rect 246528 260438 246708 260526
rect 246816 260438 246996 260526
rect 247104 260438 247284 260526
rect 247392 260438 247572 260526
rect 247680 260438 247860 260526
rect 248114 260438 248294 260526
rect 248402 260438 248582 260526
rect 248690 260438 248870 260526
rect 248978 260438 249158 260526
rect 249266 260438 249446 260526
rect 249554 260438 249734 260526
rect 249842 260438 250022 260526
rect 250130 260438 250310 260526
rect 250564 260438 250744 260526
rect 360436 260438 360560 260526
rect 360814 260438 360994 260526
rect 361102 260438 361282 260526
rect 361390 260438 361570 260526
rect 361678 260438 361858 260526
rect 361966 260438 362146 260526
rect 362254 260438 362434 260526
rect 362542 260438 362722 260526
rect 362830 260438 363010 260526
rect 363264 260438 363444 260526
rect 363552 260438 363732 260526
rect 363840 260438 364020 260526
rect 364128 260438 364308 260526
rect 364416 260438 364596 260526
rect 364704 260438 364884 260526
rect 364992 260438 365172 260526
rect 365280 260438 365460 260526
rect 365714 260438 365894 260526
rect 366002 260438 366182 260526
rect 366290 260438 366470 260526
rect 366578 260438 366758 260526
rect 366866 260438 367046 260526
rect 367154 260438 367334 260526
rect 367442 260438 367622 260526
rect 367730 260438 367910 260526
rect 243214 259962 243394 260050
rect 243502 259962 243682 260050
rect 243790 259962 243970 260050
rect 244078 259962 244258 260050
rect 244366 259962 244546 260050
rect 244654 259962 244834 260050
rect 244942 259962 245122 260050
rect 245230 259962 245410 260050
rect 245664 259962 245844 260050
rect 245952 259962 246132 260050
rect 246240 259962 246420 260050
rect 246528 259962 246708 260050
rect 246816 259962 246996 260050
rect 247104 259962 247284 260050
rect 247392 259962 247572 260050
rect 247680 259962 247860 260050
rect 248114 259962 248294 260050
rect 248402 259962 248582 260050
rect 248690 259962 248870 260050
rect 248978 259962 249158 260050
rect 249266 259962 249446 260050
rect 249554 259962 249734 260050
rect 249842 259962 250022 260050
rect 250130 259962 250310 260050
rect 250564 259962 250744 260050
rect 360436 259962 360560 260050
rect 360814 259962 360994 260050
rect 361102 259962 361282 260050
rect 361390 259962 361570 260050
rect 361678 259962 361858 260050
rect 361966 259962 362146 260050
rect 362254 259962 362434 260050
rect 362542 259962 362722 260050
rect 362830 259962 363010 260050
rect 363264 259962 363444 260050
rect 363552 259962 363732 260050
rect 363840 259962 364020 260050
rect 364128 259962 364308 260050
rect 364416 259962 364596 260050
rect 364704 259962 364884 260050
rect 364992 259962 365172 260050
rect 365280 259962 365460 260050
rect 365714 259962 365894 260050
rect 366002 259962 366182 260050
rect 366290 259962 366470 260050
rect 366578 259962 366758 260050
rect 366866 259962 367046 260050
rect 367154 259962 367334 260050
rect 367442 259962 367622 260050
rect 367730 259962 367910 260050
rect 243214 259746 243394 259834
rect 243502 259746 243682 259834
rect 243790 259746 243970 259834
rect 244078 259746 244258 259834
rect 244366 259746 244546 259834
rect 244654 259746 244834 259834
rect 244942 259746 245122 259834
rect 245230 259746 245410 259834
rect 245664 259746 245844 259834
rect 245952 259746 246132 259834
rect 246240 259746 246420 259834
rect 246528 259746 246708 259834
rect 246816 259746 246996 259834
rect 247104 259746 247284 259834
rect 247392 259746 247572 259834
rect 247680 259746 247860 259834
rect 248114 259746 248294 259834
rect 248402 259746 248582 259834
rect 248690 259746 248870 259834
rect 248978 259746 249158 259834
rect 249266 259746 249446 259834
rect 249554 259746 249734 259834
rect 249842 259746 250022 259834
rect 250130 259746 250310 259834
rect 250564 259746 250744 259834
rect 360436 259746 360560 259834
rect 360814 259746 360994 259834
rect 361102 259746 361282 259834
rect 361390 259746 361570 259834
rect 361678 259746 361858 259834
rect 361966 259746 362146 259834
rect 362254 259746 362434 259834
rect 362542 259746 362722 259834
rect 362830 259746 363010 259834
rect 363264 259746 363444 259834
rect 363552 259746 363732 259834
rect 363840 259746 364020 259834
rect 364128 259746 364308 259834
rect 364416 259746 364596 259834
rect 364704 259746 364884 259834
rect 364992 259746 365172 259834
rect 365280 259746 365460 259834
rect 365714 259746 365894 259834
rect 366002 259746 366182 259834
rect 366290 259746 366470 259834
rect 366578 259746 366758 259834
rect 366866 259746 367046 259834
rect 367154 259746 367334 259834
rect 367442 259746 367622 259834
rect 367730 259746 367910 259834
rect 243214 259270 243394 259358
rect 243502 259270 243682 259358
rect 243790 259270 243970 259358
rect 244078 259270 244258 259358
rect 244366 259270 244546 259358
rect 244654 259270 244834 259358
rect 244942 259270 245122 259358
rect 245230 259270 245410 259358
rect 245664 259270 245844 259358
rect 245952 259270 246132 259358
rect 246240 259270 246420 259358
rect 246528 259270 246708 259358
rect 246816 259270 246996 259358
rect 247104 259270 247284 259358
rect 247392 259270 247572 259358
rect 247680 259270 247860 259358
rect 248114 259270 248294 259358
rect 248402 259270 248582 259358
rect 248690 259270 248870 259358
rect 248978 259270 249158 259358
rect 249266 259270 249446 259358
rect 249554 259270 249734 259358
rect 249842 259270 250022 259358
rect 250130 259270 250310 259358
rect 250564 259270 250744 259358
rect 360436 259270 360560 259358
rect 360814 259270 360994 259358
rect 361102 259270 361282 259358
rect 361390 259270 361570 259358
rect 361678 259270 361858 259358
rect 361966 259270 362146 259358
rect 362254 259270 362434 259358
rect 362542 259270 362722 259358
rect 362830 259270 363010 259358
rect 363264 259270 363444 259358
rect 363552 259270 363732 259358
rect 363840 259270 364020 259358
rect 364128 259270 364308 259358
rect 364416 259270 364596 259358
rect 364704 259270 364884 259358
rect 364992 259270 365172 259358
rect 365280 259270 365460 259358
rect 365714 259270 365894 259358
rect 366002 259270 366182 259358
rect 366290 259270 366470 259358
rect 366578 259270 366758 259358
rect 366866 259270 367046 259358
rect 367154 259270 367334 259358
rect 367442 259270 367622 259358
rect 367730 259270 367910 259358
rect 243214 259054 243394 259142
rect 243502 259054 243682 259142
rect 243790 259054 243970 259142
rect 244078 259054 244258 259142
rect 244366 259054 244546 259142
rect 244654 259054 244834 259142
rect 244942 259054 245122 259142
rect 245230 259054 245410 259142
rect 245664 259054 245844 259142
rect 245952 259054 246132 259142
rect 246240 259054 246420 259142
rect 246528 259054 246708 259142
rect 246816 259054 246996 259142
rect 247104 259054 247284 259142
rect 247392 259054 247572 259142
rect 247680 259054 247860 259142
rect 248114 259054 248294 259142
rect 248402 259054 248582 259142
rect 248690 259054 248870 259142
rect 248978 259054 249158 259142
rect 249266 259054 249446 259142
rect 249554 259054 249734 259142
rect 249842 259054 250022 259142
rect 250130 259054 250310 259142
rect 250564 259054 250744 259142
rect 360436 259054 360560 259142
rect 360814 259054 360994 259142
rect 361102 259054 361282 259142
rect 361390 259054 361570 259142
rect 361678 259054 361858 259142
rect 361966 259054 362146 259142
rect 362254 259054 362434 259142
rect 362542 259054 362722 259142
rect 362830 259054 363010 259142
rect 363264 259054 363444 259142
rect 363552 259054 363732 259142
rect 363840 259054 364020 259142
rect 364128 259054 364308 259142
rect 364416 259054 364596 259142
rect 364704 259054 364884 259142
rect 364992 259054 365172 259142
rect 365280 259054 365460 259142
rect 365714 259054 365894 259142
rect 366002 259054 366182 259142
rect 366290 259054 366470 259142
rect 366578 259054 366758 259142
rect 366866 259054 367046 259142
rect 367154 259054 367334 259142
rect 367442 259054 367622 259142
rect 367730 259054 367910 259142
rect 243214 258578 243394 258666
rect 243502 258578 243682 258666
rect 243790 258578 243970 258666
rect 244078 258578 244258 258666
rect 244366 258578 244546 258666
rect 244654 258578 244834 258666
rect 244942 258578 245122 258666
rect 245230 258578 245410 258666
rect 245664 258578 245844 258666
rect 245952 258578 246132 258666
rect 246240 258578 246420 258666
rect 246528 258578 246708 258666
rect 246816 258578 246996 258666
rect 247104 258578 247284 258666
rect 247392 258578 247572 258666
rect 247680 258578 247860 258666
rect 248114 258578 248294 258666
rect 248402 258578 248582 258666
rect 248690 258578 248870 258666
rect 248978 258578 249158 258666
rect 249266 258578 249446 258666
rect 249554 258578 249734 258666
rect 249842 258578 250022 258666
rect 250130 258578 250310 258666
rect 250564 258578 250744 258666
rect 360436 258578 360560 258666
rect 360814 258578 360994 258666
rect 361102 258578 361282 258666
rect 361390 258578 361570 258666
rect 361678 258578 361858 258666
rect 361966 258578 362146 258666
rect 362254 258578 362434 258666
rect 362542 258578 362722 258666
rect 362830 258578 363010 258666
rect 363264 258578 363444 258666
rect 363552 258578 363732 258666
rect 363840 258578 364020 258666
rect 364128 258578 364308 258666
rect 364416 258578 364596 258666
rect 364704 258578 364884 258666
rect 364992 258578 365172 258666
rect 365280 258578 365460 258666
rect 365714 258578 365894 258666
rect 366002 258578 366182 258666
rect 366290 258578 366470 258666
rect 366578 258578 366758 258666
rect 366866 258578 367046 258666
rect 367154 258578 367334 258666
rect 367442 258578 367622 258666
rect 367730 258578 367910 258666
rect 243214 258362 243394 258450
rect 243502 258362 243682 258450
rect 243790 258362 243970 258450
rect 244078 258362 244258 258450
rect 244366 258362 244546 258450
rect 244654 258362 244834 258450
rect 244942 258362 245122 258450
rect 245230 258362 245410 258450
rect 245664 258362 245844 258450
rect 245952 258362 246132 258450
rect 246240 258362 246420 258450
rect 246528 258362 246708 258450
rect 246816 258362 246996 258450
rect 247104 258362 247284 258450
rect 247392 258362 247572 258450
rect 247680 258362 247860 258450
rect 248114 258362 248294 258450
rect 248402 258362 248582 258450
rect 248690 258362 248870 258450
rect 248978 258362 249158 258450
rect 249266 258362 249446 258450
rect 249554 258362 249734 258450
rect 249842 258362 250022 258450
rect 250130 258362 250310 258450
rect 250564 258362 250744 258450
rect 360436 258362 360560 258450
rect 360814 258362 360994 258450
rect 361102 258362 361282 258450
rect 361390 258362 361570 258450
rect 361678 258362 361858 258450
rect 361966 258362 362146 258450
rect 362254 258362 362434 258450
rect 362542 258362 362722 258450
rect 362830 258362 363010 258450
rect 363264 258362 363444 258450
rect 363552 258362 363732 258450
rect 363840 258362 364020 258450
rect 364128 258362 364308 258450
rect 364416 258362 364596 258450
rect 364704 258362 364884 258450
rect 364992 258362 365172 258450
rect 365280 258362 365460 258450
rect 365714 258362 365894 258450
rect 366002 258362 366182 258450
rect 366290 258362 366470 258450
rect 366578 258362 366758 258450
rect 366866 258362 367046 258450
rect 367154 258362 367334 258450
rect 367442 258362 367622 258450
rect 367730 258362 367910 258450
rect 243214 257886 243394 257974
rect 243502 257886 243682 257974
rect 243790 257886 243970 257974
rect 244078 257886 244258 257974
rect 244366 257886 244546 257974
rect 244654 257886 244834 257974
rect 244942 257886 245122 257974
rect 245230 257886 245410 257974
rect 245664 257886 245844 257974
rect 245952 257886 246132 257974
rect 246240 257886 246420 257974
rect 246528 257886 246708 257974
rect 246816 257886 246996 257974
rect 247104 257886 247284 257974
rect 247392 257886 247572 257974
rect 247680 257886 247860 257974
rect 248114 257886 248294 257974
rect 248402 257886 248582 257974
rect 248690 257886 248870 257974
rect 248978 257886 249158 257974
rect 249266 257886 249446 257974
rect 249554 257886 249734 257974
rect 249842 257886 250022 257974
rect 250130 257886 250310 257974
rect 250564 257886 250744 257974
rect 360436 257886 360560 257974
rect 360814 257886 360994 257974
rect 361102 257886 361282 257974
rect 361390 257886 361570 257974
rect 361678 257886 361858 257974
rect 361966 257886 362146 257974
rect 362254 257886 362434 257974
rect 362542 257886 362722 257974
rect 362830 257886 363010 257974
rect 363264 257886 363444 257974
rect 363552 257886 363732 257974
rect 363840 257886 364020 257974
rect 364128 257886 364308 257974
rect 364416 257886 364596 257974
rect 364704 257886 364884 257974
rect 364992 257886 365172 257974
rect 365280 257886 365460 257974
rect 365714 257886 365894 257974
rect 366002 257886 366182 257974
rect 366290 257886 366470 257974
rect 366578 257886 366758 257974
rect 366866 257886 367046 257974
rect 367154 257886 367334 257974
rect 367442 257886 367622 257974
rect 367730 257886 367910 257974
rect 243214 257412 243394 257500
rect 243502 257412 243682 257500
rect 243790 257412 243970 257500
rect 244078 257412 244258 257500
rect 244366 257412 244546 257500
rect 244654 257412 244834 257500
rect 244942 257412 245122 257500
rect 245230 257412 245410 257500
rect 245664 257412 245844 257500
rect 245952 257412 246132 257500
rect 246240 257412 246420 257500
rect 246528 257412 246708 257500
rect 246816 257412 246996 257500
rect 247104 257412 247284 257500
rect 247392 257412 247572 257500
rect 247680 257412 247860 257500
rect 248114 257412 248294 257500
rect 248402 257412 248582 257500
rect 248690 257412 248870 257500
rect 248978 257412 249158 257500
rect 249266 257412 249446 257500
rect 249554 257412 249734 257500
rect 249842 257412 250022 257500
rect 250130 257412 250310 257500
rect 250564 257412 250744 257500
rect 360436 257412 360560 257500
rect 360814 257412 360994 257500
rect 361102 257412 361282 257500
rect 361390 257412 361570 257500
rect 361678 257412 361858 257500
rect 361966 257412 362146 257500
rect 362254 257412 362434 257500
rect 362542 257412 362722 257500
rect 362830 257412 363010 257500
rect 363264 257412 363444 257500
rect 363552 257412 363732 257500
rect 363840 257412 364020 257500
rect 364128 257412 364308 257500
rect 364416 257412 364596 257500
rect 364704 257412 364884 257500
rect 364992 257412 365172 257500
rect 365280 257412 365460 257500
rect 365714 257412 365894 257500
rect 366002 257412 366182 257500
rect 366290 257412 366470 257500
rect 366578 257412 366758 257500
rect 366866 257412 367046 257500
rect 367154 257412 367334 257500
rect 367442 257412 367622 257500
rect 367730 257412 367910 257500
rect 243214 256936 243394 257024
rect 243502 256936 243682 257024
rect 243790 256936 243970 257024
rect 244078 256936 244258 257024
rect 244366 256936 244546 257024
rect 244654 256936 244834 257024
rect 244942 256936 245122 257024
rect 245230 256936 245410 257024
rect 245664 256936 245844 257024
rect 245952 256936 246132 257024
rect 246240 256936 246420 257024
rect 246528 256936 246708 257024
rect 246816 256936 246996 257024
rect 247104 256936 247284 257024
rect 247392 256936 247572 257024
rect 247680 256936 247860 257024
rect 248114 256936 248294 257024
rect 248402 256936 248582 257024
rect 248690 256936 248870 257024
rect 248978 256936 249158 257024
rect 249266 256936 249446 257024
rect 249554 256936 249734 257024
rect 249842 256936 250022 257024
rect 250130 256936 250310 257024
rect 250564 256936 250744 257024
rect 360436 256936 360560 257024
rect 360814 256936 360994 257024
rect 361102 256936 361282 257024
rect 361390 256936 361570 257024
rect 361678 256936 361858 257024
rect 361966 256936 362146 257024
rect 362254 256936 362434 257024
rect 362542 256936 362722 257024
rect 362830 256936 363010 257024
rect 363264 256936 363444 257024
rect 363552 256936 363732 257024
rect 363840 256936 364020 257024
rect 364128 256936 364308 257024
rect 364416 256936 364596 257024
rect 364704 256936 364884 257024
rect 364992 256936 365172 257024
rect 365280 256936 365460 257024
rect 365714 256936 365894 257024
rect 366002 256936 366182 257024
rect 366290 256936 366470 257024
rect 366578 256936 366758 257024
rect 366866 256936 367046 257024
rect 367154 256936 367334 257024
rect 367442 256936 367622 257024
rect 367730 256936 367910 257024
rect 243214 256720 243394 256808
rect 243502 256720 243682 256808
rect 243790 256720 243970 256808
rect 244078 256720 244258 256808
rect 244366 256720 244546 256808
rect 244654 256720 244834 256808
rect 244942 256720 245122 256808
rect 245230 256720 245410 256808
rect 245664 256720 245844 256808
rect 245952 256720 246132 256808
rect 246240 256720 246420 256808
rect 246528 256720 246708 256808
rect 246816 256720 246996 256808
rect 247104 256720 247284 256808
rect 247392 256720 247572 256808
rect 247680 256720 247860 256808
rect 248114 256720 248294 256808
rect 248402 256720 248582 256808
rect 248690 256720 248870 256808
rect 248978 256720 249158 256808
rect 249266 256720 249446 256808
rect 249554 256720 249734 256808
rect 249842 256720 250022 256808
rect 250130 256720 250310 256808
rect 250564 256720 250744 256808
rect 360436 256720 360560 256808
rect 360814 256720 360994 256808
rect 361102 256720 361282 256808
rect 361390 256720 361570 256808
rect 361678 256720 361858 256808
rect 361966 256720 362146 256808
rect 362254 256720 362434 256808
rect 362542 256720 362722 256808
rect 362830 256720 363010 256808
rect 363264 256720 363444 256808
rect 363552 256720 363732 256808
rect 363840 256720 364020 256808
rect 364128 256720 364308 256808
rect 364416 256720 364596 256808
rect 364704 256720 364884 256808
rect 364992 256720 365172 256808
rect 365280 256720 365460 256808
rect 365714 256720 365894 256808
rect 366002 256720 366182 256808
rect 366290 256720 366470 256808
rect 366578 256720 366758 256808
rect 366866 256720 367046 256808
rect 367154 256720 367334 256808
rect 367442 256720 367622 256808
rect 367730 256720 367910 256808
rect 243214 256244 243394 256332
rect 243502 256244 243682 256332
rect 243790 256244 243970 256332
rect 244078 256244 244258 256332
rect 244366 256244 244546 256332
rect 244654 256244 244834 256332
rect 244942 256244 245122 256332
rect 245230 256244 245410 256332
rect 245664 256244 245844 256332
rect 245952 256244 246132 256332
rect 246240 256244 246420 256332
rect 246528 256244 246708 256332
rect 246816 256244 246996 256332
rect 247104 256244 247284 256332
rect 247392 256244 247572 256332
rect 247680 256244 247860 256332
rect 248114 256244 248294 256332
rect 248402 256244 248582 256332
rect 248690 256244 248870 256332
rect 248978 256244 249158 256332
rect 249266 256244 249446 256332
rect 249554 256244 249734 256332
rect 249842 256244 250022 256332
rect 250130 256244 250310 256332
rect 250564 256244 250744 256332
rect 360436 256244 360560 256332
rect 360814 256244 360994 256332
rect 361102 256244 361282 256332
rect 361390 256244 361570 256332
rect 361678 256244 361858 256332
rect 361966 256244 362146 256332
rect 362254 256244 362434 256332
rect 362542 256244 362722 256332
rect 362830 256244 363010 256332
rect 363264 256244 363444 256332
rect 363552 256244 363732 256332
rect 363840 256244 364020 256332
rect 364128 256244 364308 256332
rect 364416 256244 364596 256332
rect 364704 256244 364884 256332
rect 364992 256244 365172 256332
rect 365280 256244 365460 256332
rect 365714 256244 365894 256332
rect 366002 256244 366182 256332
rect 366290 256244 366470 256332
rect 366578 256244 366758 256332
rect 366866 256244 367046 256332
rect 367154 256244 367334 256332
rect 367442 256244 367622 256332
rect 367730 256244 367910 256332
rect 243214 256028 243394 256116
rect 243502 256028 243682 256116
rect 243790 256028 243970 256116
rect 244078 256028 244258 256116
rect 244366 256028 244546 256116
rect 244654 256028 244834 256116
rect 244942 256028 245122 256116
rect 245230 256028 245410 256116
rect 245664 256028 245844 256116
rect 245952 256028 246132 256116
rect 246240 256028 246420 256116
rect 246528 256028 246708 256116
rect 246816 256028 246996 256116
rect 247104 256028 247284 256116
rect 247392 256028 247572 256116
rect 247680 256028 247860 256116
rect 248114 256028 248294 256116
rect 248402 256028 248582 256116
rect 248690 256028 248870 256116
rect 248978 256028 249158 256116
rect 249266 256028 249446 256116
rect 249554 256028 249734 256116
rect 249842 256028 250022 256116
rect 250130 256028 250310 256116
rect 250564 256028 250744 256116
rect 360436 256028 360560 256116
rect 360814 256028 360994 256116
rect 361102 256028 361282 256116
rect 361390 256028 361570 256116
rect 361678 256028 361858 256116
rect 361966 256028 362146 256116
rect 362254 256028 362434 256116
rect 362542 256028 362722 256116
rect 362830 256028 363010 256116
rect 363264 256028 363444 256116
rect 363552 256028 363732 256116
rect 363840 256028 364020 256116
rect 364128 256028 364308 256116
rect 364416 256028 364596 256116
rect 364704 256028 364884 256116
rect 364992 256028 365172 256116
rect 365280 256028 365460 256116
rect 365714 256028 365894 256116
rect 366002 256028 366182 256116
rect 366290 256028 366470 256116
rect 366578 256028 366758 256116
rect 366866 256028 367046 256116
rect 367154 256028 367334 256116
rect 367442 256028 367622 256116
rect 367730 256028 367910 256116
rect 243214 255552 243394 255640
rect 243502 255552 243682 255640
rect 243790 255552 243970 255640
rect 244078 255552 244258 255640
rect 244366 255552 244546 255640
rect 244654 255552 244834 255640
rect 244942 255552 245122 255640
rect 245230 255552 245410 255640
rect 245664 255552 245844 255640
rect 245952 255552 246132 255640
rect 246240 255552 246420 255640
rect 246528 255552 246708 255640
rect 246816 255552 246996 255640
rect 247104 255552 247284 255640
rect 247392 255552 247572 255640
rect 247680 255552 247860 255640
rect 248114 255552 248294 255640
rect 248402 255552 248582 255640
rect 248690 255552 248870 255640
rect 248978 255552 249158 255640
rect 249266 255552 249446 255640
rect 249554 255552 249734 255640
rect 249842 255552 250022 255640
rect 250130 255552 250310 255640
rect 250564 255552 250744 255640
rect 360436 255552 360560 255640
rect 360814 255552 360994 255640
rect 361102 255552 361282 255640
rect 361390 255552 361570 255640
rect 361678 255552 361858 255640
rect 361966 255552 362146 255640
rect 362254 255552 362434 255640
rect 362542 255552 362722 255640
rect 362830 255552 363010 255640
rect 363264 255552 363444 255640
rect 363552 255552 363732 255640
rect 363840 255552 364020 255640
rect 364128 255552 364308 255640
rect 364416 255552 364596 255640
rect 364704 255552 364884 255640
rect 364992 255552 365172 255640
rect 365280 255552 365460 255640
rect 365714 255552 365894 255640
rect 366002 255552 366182 255640
rect 366290 255552 366470 255640
rect 366578 255552 366758 255640
rect 366866 255552 367046 255640
rect 367154 255552 367334 255640
rect 367442 255552 367622 255640
rect 367730 255552 367910 255640
rect 243214 255336 243394 255424
rect 243502 255336 243682 255424
rect 243790 255336 243970 255424
rect 244078 255336 244258 255424
rect 244366 255336 244546 255424
rect 244654 255336 244834 255424
rect 244942 255336 245122 255424
rect 245230 255336 245410 255424
rect 245664 255336 245844 255424
rect 245952 255336 246132 255424
rect 246240 255336 246420 255424
rect 246528 255336 246708 255424
rect 246816 255336 246996 255424
rect 247104 255336 247284 255424
rect 247392 255336 247572 255424
rect 247680 255336 247860 255424
rect 248114 255336 248294 255424
rect 248402 255336 248582 255424
rect 248690 255336 248870 255424
rect 248978 255336 249158 255424
rect 249266 255336 249446 255424
rect 249554 255336 249734 255424
rect 249842 255336 250022 255424
rect 250130 255336 250310 255424
rect 250564 255336 250744 255424
rect 360436 255336 360560 255424
rect 360814 255336 360994 255424
rect 361102 255336 361282 255424
rect 361390 255336 361570 255424
rect 361678 255336 361858 255424
rect 361966 255336 362146 255424
rect 362254 255336 362434 255424
rect 362542 255336 362722 255424
rect 362830 255336 363010 255424
rect 363264 255336 363444 255424
rect 363552 255336 363732 255424
rect 363840 255336 364020 255424
rect 364128 255336 364308 255424
rect 364416 255336 364596 255424
rect 364704 255336 364884 255424
rect 364992 255336 365172 255424
rect 365280 255336 365460 255424
rect 365714 255336 365894 255424
rect 366002 255336 366182 255424
rect 366290 255336 366470 255424
rect 366578 255336 366758 255424
rect 366866 255336 367046 255424
rect 367154 255336 367334 255424
rect 367442 255336 367622 255424
rect 367730 255336 367910 255424
rect 243214 254860 243394 254948
rect 243502 254860 243682 254948
rect 243790 254860 243970 254948
rect 244078 254860 244258 254948
rect 244366 254860 244546 254948
rect 244654 254860 244834 254948
rect 244942 254860 245122 254948
rect 245230 254860 245410 254948
rect 245664 254860 245844 254948
rect 245952 254860 246132 254948
rect 246240 254860 246420 254948
rect 246528 254860 246708 254948
rect 246816 254860 246996 254948
rect 247104 254860 247284 254948
rect 247392 254860 247572 254948
rect 247680 254860 247860 254948
rect 248114 254860 248294 254948
rect 248402 254860 248582 254948
rect 248690 254860 248870 254948
rect 248978 254860 249158 254948
rect 249266 254860 249446 254948
rect 249554 254860 249734 254948
rect 249842 254860 250022 254948
rect 250130 254860 250310 254948
rect 250564 254860 250744 254948
rect 360436 254860 360560 254948
rect 360814 254860 360994 254948
rect 361102 254860 361282 254948
rect 361390 254860 361570 254948
rect 361678 254860 361858 254948
rect 361966 254860 362146 254948
rect 362254 254860 362434 254948
rect 362542 254860 362722 254948
rect 362830 254860 363010 254948
rect 363264 254860 363444 254948
rect 363552 254860 363732 254948
rect 363840 254860 364020 254948
rect 364128 254860 364308 254948
rect 364416 254860 364596 254948
rect 364704 254860 364884 254948
rect 364992 254860 365172 254948
rect 365280 254860 365460 254948
rect 365714 254860 365894 254948
rect 366002 254860 366182 254948
rect 366290 254860 366470 254948
rect 366578 254860 366758 254948
rect 366866 254860 367046 254948
rect 367154 254860 367334 254948
rect 367442 254860 367622 254948
rect 367730 254860 367910 254948
rect 243214 254386 243394 254474
rect 243502 254386 243682 254474
rect 243790 254386 243970 254474
rect 244078 254386 244258 254474
rect 244366 254386 244546 254474
rect 244654 254386 244834 254474
rect 244942 254386 245122 254474
rect 245230 254386 245410 254474
rect 245664 254386 245844 254474
rect 245952 254386 246132 254474
rect 246240 254386 246420 254474
rect 246528 254386 246708 254474
rect 246816 254386 246996 254474
rect 247104 254386 247284 254474
rect 247392 254386 247572 254474
rect 247680 254386 247860 254474
rect 248114 254386 248294 254474
rect 248402 254386 248582 254474
rect 248690 254386 248870 254474
rect 248978 254386 249158 254474
rect 249266 254386 249446 254474
rect 249554 254386 249734 254474
rect 249842 254386 250022 254474
rect 250130 254386 250310 254474
rect 250564 254386 250744 254474
rect 360436 254386 360560 254474
rect 360814 254386 360994 254474
rect 361102 254386 361282 254474
rect 361390 254386 361570 254474
rect 361678 254386 361858 254474
rect 361966 254386 362146 254474
rect 362254 254386 362434 254474
rect 362542 254386 362722 254474
rect 362830 254386 363010 254474
rect 363264 254386 363444 254474
rect 363552 254386 363732 254474
rect 363840 254386 364020 254474
rect 364128 254386 364308 254474
rect 364416 254386 364596 254474
rect 364704 254386 364884 254474
rect 364992 254386 365172 254474
rect 365280 254386 365460 254474
rect 365714 254386 365894 254474
rect 366002 254386 366182 254474
rect 366290 254386 366470 254474
rect 366578 254386 366758 254474
rect 366866 254386 367046 254474
rect 367154 254386 367334 254474
rect 367442 254386 367622 254474
rect 367730 254386 367910 254474
rect 243214 253910 243394 253998
rect 243502 253910 243682 253998
rect 243790 253910 243970 253998
rect 244078 253910 244258 253998
rect 244366 253910 244546 253998
rect 244654 253910 244834 253998
rect 244942 253910 245122 253998
rect 245230 253910 245410 253998
rect 245664 253910 245844 253998
rect 245952 253910 246132 253998
rect 246240 253910 246420 253998
rect 246528 253910 246708 253998
rect 246816 253910 246996 253998
rect 247104 253910 247284 253998
rect 247392 253910 247572 253998
rect 247680 253910 247860 253998
rect 248114 253910 248294 253998
rect 248402 253910 248582 253998
rect 248690 253910 248870 253998
rect 248978 253910 249158 253998
rect 249266 253910 249446 253998
rect 249554 253910 249734 253998
rect 249842 253910 250022 253998
rect 250130 253910 250310 253998
rect 250564 253910 250744 253998
rect 360436 253910 360560 253998
rect 360814 253910 360994 253998
rect 361102 253910 361282 253998
rect 361390 253910 361570 253998
rect 361678 253910 361858 253998
rect 361966 253910 362146 253998
rect 362254 253910 362434 253998
rect 362542 253910 362722 253998
rect 362830 253910 363010 253998
rect 363264 253910 363444 253998
rect 363552 253910 363732 253998
rect 363840 253910 364020 253998
rect 364128 253910 364308 253998
rect 364416 253910 364596 253998
rect 364704 253910 364884 253998
rect 364992 253910 365172 253998
rect 365280 253910 365460 253998
rect 365714 253910 365894 253998
rect 366002 253910 366182 253998
rect 366290 253910 366470 253998
rect 366578 253910 366758 253998
rect 366866 253910 367046 253998
rect 367154 253910 367334 253998
rect 367442 253910 367622 253998
rect 367730 253910 367910 253998
rect 243214 253694 243394 253782
rect 243502 253694 243682 253782
rect 243790 253694 243970 253782
rect 244078 253694 244258 253782
rect 244366 253694 244546 253782
rect 244654 253694 244834 253782
rect 244942 253694 245122 253782
rect 245230 253694 245410 253782
rect 245664 253694 245844 253782
rect 245952 253694 246132 253782
rect 246240 253694 246420 253782
rect 246528 253694 246708 253782
rect 246816 253694 246996 253782
rect 247104 253694 247284 253782
rect 247392 253694 247572 253782
rect 247680 253694 247860 253782
rect 248114 253694 248294 253782
rect 248402 253694 248582 253782
rect 248690 253694 248870 253782
rect 248978 253694 249158 253782
rect 249266 253694 249446 253782
rect 249554 253694 249734 253782
rect 249842 253694 250022 253782
rect 250130 253694 250310 253782
rect 250564 253694 250744 253782
rect 360436 253694 360560 253782
rect 360814 253694 360994 253782
rect 361102 253694 361282 253782
rect 361390 253694 361570 253782
rect 361678 253694 361858 253782
rect 361966 253694 362146 253782
rect 362254 253694 362434 253782
rect 362542 253694 362722 253782
rect 362830 253694 363010 253782
rect 363264 253694 363444 253782
rect 363552 253694 363732 253782
rect 363840 253694 364020 253782
rect 364128 253694 364308 253782
rect 364416 253694 364596 253782
rect 364704 253694 364884 253782
rect 364992 253694 365172 253782
rect 365280 253694 365460 253782
rect 365714 253694 365894 253782
rect 366002 253694 366182 253782
rect 366290 253694 366470 253782
rect 366578 253694 366758 253782
rect 366866 253694 367046 253782
rect 367154 253694 367334 253782
rect 367442 253694 367622 253782
rect 367730 253694 367910 253782
rect 243214 253218 243394 253306
rect 243502 253218 243682 253306
rect 243790 253218 243970 253306
rect 244078 253218 244258 253306
rect 244366 253218 244546 253306
rect 244654 253218 244834 253306
rect 244942 253218 245122 253306
rect 245230 253218 245410 253306
rect 245664 253218 245844 253306
rect 245952 253218 246132 253306
rect 246240 253218 246420 253306
rect 246528 253218 246708 253306
rect 246816 253218 246996 253306
rect 247104 253218 247284 253306
rect 247392 253218 247572 253306
rect 247680 253218 247860 253306
rect 248114 253218 248294 253306
rect 248402 253218 248582 253306
rect 248690 253218 248870 253306
rect 248978 253218 249158 253306
rect 249266 253218 249446 253306
rect 249554 253218 249734 253306
rect 249842 253218 250022 253306
rect 250130 253218 250310 253306
rect 250564 253218 250744 253306
rect 360436 253218 360560 253306
rect 360814 253218 360994 253306
rect 361102 253218 361282 253306
rect 361390 253218 361570 253306
rect 361678 253218 361858 253306
rect 361966 253218 362146 253306
rect 362254 253218 362434 253306
rect 362542 253218 362722 253306
rect 362830 253218 363010 253306
rect 363264 253218 363444 253306
rect 363552 253218 363732 253306
rect 363840 253218 364020 253306
rect 364128 253218 364308 253306
rect 364416 253218 364596 253306
rect 364704 253218 364884 253306
rect 364992 253218 365172 253306
rect 365280 253218 365460 253306
rect 365714 253218 365894 253306
rect 366002 253218 366182 253306
rect 366290 253218 366470 253306
rect 366578 253218 366758 253306
rect 366866 253218 367046 253306
rect 367154 253218 367334 253306
rect 367442 253218 367622 253306
rect 367730 253218 367910 253306
rect 243214 253002 243394 253090
rect 243502 253002 243682 253090
rect 243790 253002 243970 253090
rect 244078 253002 244258 253090
rect 244366 253002 244546 253090
rect 244654 253002 244834 253090
rect 244942 253002 245122 253090
rect 245230 253002 245410 253090
rect 245664 253002 245844 253090
rect 245952 253002 246132 253090
rect 246240 253002 246420 253090
rect 246528 253002 246708 253090
rect 246816 253002 246996 253090
rect 247104 253002 247284 253090
rect 247392 253002 247572 253090
rect 247680 253002 247860 253090
rect 248114 253002 248294 253090
rect 248402 253002 248582 253090
rect 248690 253002 248870 253090
rect 248978 253002 249158 253090
rect 249266 253002 249446 253090
rect 249554 253002 249734 253090
rect 249842 253002 250022 253090
rect 250130 253002 250310 253090
rect 250564 253002 250744 253090
rect 360436 253002 360560 253090
rect 360814 253002 360994 253090
rect 361102 253002 361282 253090
rect 361390 253002 361570 253090
rect 361678 253002 361858 253090
rect 361966 253002 362146 253090
rect 362254 253002 362434 253090
rect 362542 253002 362722 253090
rect 362830 253002 363010 253090
rect 363264 253002 363444 253090
rect 363552 253002 363732 253090
rect 363840 253002 364020 253090
rect 364128 253002 364308 253090
rect 364416 253002 364596 253090
rect 364704 253002 364884 253090
rect 364992 253002 365172 253090
rect 365280 253002 365460 253090
rect 365714 253002 365894 253090
rect 366002 253002 366182 253090
rect 366290 253002 366470 253090
rect 366578 253002 366758 253090
rect 366866 253002 367046 253090
rect 367154 253002 367334 253090
rect 367442 253002 367622 253090
rect 367730 253002 367910 253090
rect 243214 252526 243394 252614
rect 243502 252526 243682 252614
rect 243790 252526 243970 252614
rect 244078 252526 244258 252614
rect 244366 252526 244546 252614
rect 244654 252526 244834 252614
rect 244942 252526 245122 252614
rect 245230 252526 245410 252614
rect 245664 252526 245844 252614
rect 245952 252526 246132 252614
rect 246240 252526 246420 252614
rect 246528 252526 246708 252614
rect 246816 252526 246996 252614
rect 247104 252526 247284 252614
rect 247392 252526 247572 252614
rect 247680 252526 247860 252614
rect 248114 252526 248294 252614
rect 248402 252526 248582 252614
rect 248690 252526 248870 252614
rect 248978 252526 249158 252614
rect 249266 252526 249446 252614
rect 249554 252526 249734 252614
rect 249842 252526 250022 252614
rect 250130 252526 250310 252614
rect 250564 252526 250744 252614
rect 360436 252526 360560 252614
rect 360814 252526 360994 252614
rect 361102 252526 361282 252614
rect 361390 252526 361570 252614
rect 361678 252526 361858 252614
rect 361966 252526 362146 252614
rect 362254 252526 362434 252614
rect 362542 252526 362722 252614
rect 362830 252526 363010 252614
rect 363264 252526 363444 252614
rect 363552 252526 363732 252614
rect 363840 252526 364020 252614
rect 364128 252526 364308 252614
rect 364416 252526 364596 252614
rect 364704 252526 364884 252614
rect 364992 252526 365172 252614
rect 365280 252526 365460 252614
rect 365714 252526 365894 252614
rect 366002 252526 366182 252614
rect 366290 252526 366470 252614
rect 366578 252526 366758 252614
rect 366866 252526 367046 252614
rect 367154 252526 367334 252614
rect 367442 252526 367622 252614
rect 367730 252526 367910 252614
rect 243214 252310 243394 252398
rect 243502 252310 243682 252398
rect 243790 252310 243970 252398
rect 244078 252310 244258 252398
rect 244366 252310 244546 252398
rect 244654 252310 244834 252398
rect 244942 252310 245122 252398
rect 245230 252310 245410 252398
rect 245664 252310 245844 252398
rect 245952 252310 246132 252398
rect 246240 252310 246420 252398
rect 246528 252310 246708 252398
rect 246816 252310 246996 252398
rect 247104 252310 247284 252398
rect 247392 252310 247572 252398
rect 247680 252310 247860 252398
rect 248114 252310 248294 252398
rect 248402 252310 248582 252398
rect 248690 252310 248870 252398
rect 248978 252310 249158 252398
rect 249266 252310 249446 252398
rect 249554 252310 249734 252398
rect 249842 252310 250022 252398
rect 250130 252310 250310 252398
rect 250564 252310 250744 252398
rect 360436 252310 360560 252398
rect 360814 252310 360994 252398
rect 361102 252310 361282 252398
rect 361390 252310 361570 252398
rect 361678 252310 361858 252398
rect 361966 252310 362146 252398
rect 362254 252310 362434 252398
rect 362542 252310 362722 252398
rect 362830 252310 363010 252398
rect 363264 252310 363444 252398
rect 363552 252310 363732 252398
rect 363840 252310 364020 252398
rect 364128 252310 364308 252398
rect 364416 252310 364596 252398
rect 364704 252310 364884 252398
rect 364992 252310 365172 252398
rect 365280 252310 365460 252398
rect 365714 252310 365894 252398
rect 366002 252310 366182 252398
rect 366290 252310 366470 252398
rect 366578 252310 366758 252398
rect 366866 252310 367046 252398
rect 367154 252310 367334 252398
rect 367442 252310 367622 252398
rect 367730 252310 367910 252398
rect 243214 251834 243394 251922
rect 243502 251834 243682 251922
rect 243790 251834 243970 251922
rect 244078 251834 244258 251922
rect 244366 251834 244546 251922
rect 244654 251834 244834 251922
rect 244942 251834 245122 251922
rect 245230 251834 245410 251922
rect 245664 251834 245844 251922
rect 245952 251834 246132 251922
rect 246240 251834 246420 251922
rect 246528 251834 246708 251922
rect 246816 251834 246996 251922
rect 247104 251834 247284 251922
rect 247392 251834 247572 251922
rect 247680 251834 247860 251922
rect 248114 251834 248294 251922
rect 248402 251834 248582 251922
rect 248690 251834 248870 251922
rect 248978 251834 249158 251922
rect 249266 251834 249446 251922
rect 249554 251834 249734 251922
rect 249842 251834 250022 251922
rect 250130 251834 250310 251922
rect 250564 251834 250744 251922
rect 360436 251834 360560 251922
rect 360814 251834 360994 251922
rect 361102 251834 361282 251922
rect 361390 251834 361570 251922
rect 361678 251834 361858 251922
rect 361966 251834 362146 251922
rect 362254 251834 362434 251922
rect 362542 251834 362722 251922
rect 362830 251834 363010 251922
rect 363264 251834 363444 251922
rect 363552 251834 363732 251922
rect 363840 251834 364020 251922
rect 364128 251834 364308 251922
rect 364416 251834 364596 251922
rect 364704 251834 364884 251922
rect 364992 251834 365172 251922
rect 365280 251834 365460 251922
rect 365714 251834 365894 251922
rect 366002 251834 366182 251922
rect 366290 251834 366470 251922
rect 366578 251834 366758 251922
rect 366866 251834 367046 251922
rect 367154 251834 367334 251922
rect 367442 251834 367622 251922
rect 367730 251834 367910 251922
rect 243214 251360 243394 251448
rect 243502 251360 243682 251448
rect 243790 251360 243970 251448
rect 244078 251360 244258 251448
rect 244366 251360 244546 251448
rect 244654 251360 244834 251448
rect 244942 251360 245122 251448
rect 245230 251360 245410 251448
rect 245664 251360 245844 251448
rect 245952 251360 246132 251448
rect 246240 251360 246420 251448
rect 246528 251360 246708 251448
rect 246816 251360 246996 251448
rect 247104 251360 247284 251448
rect 247392 251360 247572 251448
rect 247680 251360 247860 251448
rect 248114 251360 248294 251448
rect 248402 251360 248582 251448
rect 248690 251360 248870 251448
rect 248978 251360 249158 251448
rect 249266 251360 249446 251448
rect 249554 251360 249734 251448
rect 249842 251360 250022 251448
rect 250130 251360 250310 251448
rect 250564 251360 250744 251448
rect 360436 251360 360560 251448
rect 360814 251360 360994 251448
rect 361102 251360 361282 251448
rect 361390 251360 361570 251448
rect 361678 251360 361858 251448
rect 361966 251360 362146 251448
rect 362254 251360 362434 251448
rect 362542 251360 362722 251448
rect 362830 251360 363010 251448
rect 363264 251360 363444 251448
rect 363552 251360 363732 251448
rect 363840 251360 364020 251448
rect 364128 251360 364308 251448
rect 364416 251360 364596 251448
rect 364704 251360 364884 251448
rect 364992 251360 365172 251448
rect 365280 251360 365460 251448
rect 365714 251360 365894 251448
rect 366002 251360 366182 251448
rect 366290 251360 366470 251448
rect 366578 251360 366758 251448
rect 366866 251360 367046 251448
rect 367154 251360 367334 251448
rect 367442 251360 367622 251448
rect 367730 251360 367910 251448
rect 243214 250884 243394 250972
rect 243502 250884 243682 250972
rect 243790 250884 243970 250972
rect 244078 250884 244258 250972
rect 244366 250884 244546 250972
rect 244654 250884 244834 250972
rect 244942 250884 245122 250972
rect 245230 250884 245410 250972
rect 245664 250884 245844 250972
rect 245952 250884 246132 250972
rect 246240 250884 246420 250972
rect 246528 250884 246708 250972
rect 246816 250884 246996 250972
rect 247104 250884 247284 250972
rect 247392 250884 247572 250972
rect 247680 250884 247860 250972
rect 248114 250884 248294 250972
rect 248402 250884 248582 250972
rect 248690 250884 248870 250972
rect 248978 250884 249158 250972
rect 249266 250884 249446 250972
rect 249554 250884 249734 250972
rect 249842 250884 250022 250972
rect 250130 250884 250310 250972
rect 250564 250884 250744 250972
rect 360436 250884 360560 250972
rect 360814 250884 360994 250972
rect 361102 250884 361282 250972
rect 361390 250884 361570 250972
rect 361678 250884 361858 250972
rect 361966 250884 362146 250972
rect 362254 250884 362434 250972
rect 362542 250884 362722 250972
rect 362830 250884 363010 250972
rect 363264 250884 363444 250972
rect 363552 250884 363732 250972
rect 363840 250884 364020 250972
rect 364128 250884 364308 250972
rect 364416 250884 364596 250972
rect 364704 250884 364884 250972
rect 364992 250884 365172 250972
rect 365280 250884 365460 250972
rect 365714 250884 365894 250972
rect 366002 250884 366182 250972
rect 366290 250884 366470 250972
rect 366578 250884 366758 250972
rect 366866 250884 367046 250972
rect 367154 250884 367334 250972
rect 367442 250884 367622 250972
rect 367730 250884 367910 250972
rect 243214 250668 243394 250756
rect 243502 250668 243682 250756
rect 243790 250668 243970 250756
rect 244078 250668 244258 250756
rect 244366 250668 244546 250756
rect 244654 250668 244834 250756
rect 244942 250668 245122 250756
rect 245230 250668 245410 250756
rect 245664 250668 245844 250756
rect 245952 250668 246132 250756
rect 246240 250668 246420 250756
rect 246528 250668 246708 250756
rect 246816 250668 246996 250756
rect 247104 250668 247284 250756
rect 247392 250668 247572 250756
rect 247680 250668 247860 250756
rect 248114 250668 248294 250756
rect 248402 250668 248582 250756
rect 248690 250668 248870 250756
rect 248978 250668 249158 250756
rect 249266 250668 249446 250756
rect 249554 250668 249734 250756
rect 249842 250668 250022 250756
rect 250130 250668 250310 250756
rect 250564 250668 250744 250756
rect 360436 250668 360560 250756
rect 360814 250668 360994 250756
rect 361102 250668 361282 250756
rect 361390 250668 361570 250756
rect 361678 250668 361858 250756
rect 361966 250668 362146 250756
rect 362254 250668 362434 250756
rect 362542 250668 362722 250756
rect 362830 250668 363010 250756
rect 363264 250668 363444 250756
rect 363552 250668 363732 250756
rect 363840 250668 364020 250756
rect 364128 250668 364308 250756
rect 364416 250668 364596 250756
rect 364704 250668 364884 250756
rect 364992 250668 365172 250756
rect 365280 250668 365460 250756
rect 365714 250668 365894 250756
rect 366002 250668 366182 250756
rect 366290 250668 366470 250756
rect 366578 250668 366758 250756
rect 366866 250668 367046 250756
rect 367154 250668 367334 250756
rect 367442 250668 367622 250756
rect 367730 250668 367910 250756
rect 243214 250192 243394 250280
rect 243502 250192 243682 250280
rect 243790 250192 243970 250280
rect 244078 250192 244258 250280
rect 244366 250192 244546 250280
rect 244654 250192 244834 250280
rect 244942 250192 245122 250280
rect 245230 250192 245410 250280
rect 245664 250192 245844 250280
rect 245952 250192 246132 250280
rect 246240 250192 246420 250280
rect 246528 250192 246708 250280
rect 246816 250192 246996 250280
rect 247104 250192 247284 250280
rect 247392 250192 247572 250280
rect 247680 250192 247860 250280
rect 248114 250192 248294 250280
rect 248402 250192 248582 250280
rect 248690 250192 248870 250280
rect 248978 250192 249158 250280
rect 249266 250192 249446 250280
rect 249554 250192 249734 250280
rect 249842 250192 250022 250280
rect 250130 250192 250310 250280
rect 250564 250192 250744 250280
rect 360436 250192 360560 250280
rect 360814 250192 360994 250280
rect 361102 250192 361282 250280
rect 361390 250192 361570 250280
rect 361678 250192 361858 250280
rect 361966 250192 362146 250280
rect 362254 250192 362434 250280
rect 362542 250192 362722 250280
rect 362830 250192 363010 250280
rect 363264 250192 363444 250280
rect 363552 250192 363732 250280
rect 363840 250192 364020 250280
rect 364128 250192 364308 250280
rect 364416 250192 364596 250280
rect 364704 250192 364884 250280
rect 364992 250192 365172 250280
rect 365280 250192 365460 250280
rect 365714 250192 365894 250280
rect 366002 250192 366182 250280
rect 366290 250192 366470 250280
rect 366578 250192 366758 250280
rect 366866 250192 367046 250280
rect 367154 250192 367334 250280
rect 367442 250192 367622 250280
rect 367730 250192 367910 250280
rect 243214 249976 243394 250064
rect 243502 249976 243682 250064
rect 243790 249976 243970 250064
rect 244078 249976 244258 250064
rect 244366 249976 244546 250064
rect 244654 249976 244834 250064
rect 244942 249976 245122 250064
rect 245230 249976 245410 250064
rect 245664 249976 245844 250064
rect 245952 249976 246132 250064
rect 246240 249976 246420 250064
rect 246528 249976 246708 250064
rect 246816 249976 246996 250064
rect 247104 249976 247284 250064
rect 247392 249976 247572 250064
rect 247680 249976 247860 250064
rect 248114 249976 248294 250064
rect 248402 249976 248582 250064
rect 248690 249976 248870 250064
rect 248978 249976 249158 250064
rect 249266 249976 249446 250064
rect 249554 249976 249734 250064
rect 249842 249976 250022 250064
rect 250130 249976 250310 250064
rect 250564 249976 250744 250064
rect 360436 249976 360560 250064
rect 360814 249976 360994 250064
rect 361102 249976 361282 250064
rect 361390 249976 361570 250064
rect 361678 249976 361858 250064
rect 361966 249976 362146 250064
rect 362254 249976 362434 250064
rect 362542 249976 362722 250064
rect 362830 249976 363010 250064
rect 363264 249976 363444 250064
rect 363552 249976 363732 250064
rect 363840 249976 364020 250064
rect 364128 249976 364308 250064
rect 364416 249976 364596 250064
rect 364704 249976 364884 250064
rect 364992 249976 365172 250064
rect 365280 249976 365460 250064
rect 365714 249976 365894 250064
rect 366002 249976 366182 250064
rect 366290 249976 366470 250064
rect 366578 249976 366758 250064
rect 366866 249976 367046 250064
rect 367154 249976 367334 250064
rect 367442 249976 367622 250064
rect 367730 249976 367910 250064
rect 243214 249500 243394 249588
rect 243502 249500 243682 249588
rect 243790 249500 243970 249588
rect 244078 249500 244258 249588
rect 244366 249500 244546 249588
rect 244654 249500 244834 249588
rect 244942 249500 245122 249588
rect 245230 249500 245410 249588
rect 245664 249500 245844 249588
rect 245952 249500 246132 249588
rect 246240 249500 246420 249588
rect 246528 249500 246708 249588
rect 246816 249500 246996 249588
rect 247104 249500 247284 249588
rect 247392 249500 247572 249588
rect 247680 249500 247860 249588
rect 248114 249500 248294 249588
rect 248402 249500 248582 249588
rect 248690 249500 248870 249588
rect 248978 249500 249158 249588
rect 249266 249500 249446 249588
rect 249554 249500 249734 249588
rect 249842 249500 250022 249588
rect 250130 249500 250310 249588
rect 250564 249500 250744 249588
rect 360436 249500 360560 249588
rect 360814 249500 360994 249588
rect 361102 249500 361282 249588
rect 361390 249500 361570 249588
rect 361678 249500 361858 249588
rect 361966 249500 362146 249588
rect 362254 249500 362434 249588
rect 362542 249500 362722 249588
rect 362830 249500 363010 249588
rect 363264 249500 363444 249588
rect 363552 249500 363732 249588
rect 363840 249500 364020 249588
rect 364128 249500 364308 249588
rect 364416 249500 364596 249588
rect 364704 249500 364884 249588
rect 364992 249500 365172 249588
rect 365280 249500 365460 249588
rect 365714 249500 365894 249588
rect 366002 249500 366182 249588
rect 366290 249500 366470 249588
rect 366578 249500 366758 249588
rect 366866 249500 367046 249588
rect 367154 249500 367334 249588
rect 367442 249500 367622 249588
rect 367730 249500 367910 249588
rect 243214 249284 243394 249372
rect 243502 249284 243682 249372
rect 243790 249284 243970 249372
rect 244078 249284 244258 249372
rect 244366 249284 244546 249372
rect 244654 249284 244834 249372
rect 244942 249284 245122 249372
rect 245230 249284 245410 249372
rect 245664 249284 245844 249372
rect 245952 249284 246132 249372
rect 246240 249284 246420 249372
rect 246528 249284 246708 249372
rect 246816 249284 246996 249372
rect 247104 249284 247284 249372
rect 247392 249284 247572 249372
rect 247680 249284 247860 249372
rect 248114 249284 248294 249372
rect 248402 249284 248582 249372
rect 248690 249284 248870 249372
rect 248978 249284 249158 249372
rect 249266 249284 249446 249372
rect 249554 249284 249734 249372
rect 249842 249284 250022 249372
rect 250130 249284 250310 249372
rect 250564 249284 250744 249372
rect 360436 249284 360560 249372
rect 360814 249284 360994 249372
rect 361102 249284 361282 249372
rect 361390 249284 361570 249372
rect 361678 249284 361858 249372
rect 361966 249284 362146 249372
rect 362254 249284 362434 249372
rect 362542 249284 362722 249372
rect 362830 249284 363010 249372
rect 363264 249284 363444 249372
rect 363552 249284 363732 249372
rect 363840 249284 364020 249372
rect 364128 249284 364308 249372
rect 364416 249284 364596 249372
rect 364704 249284 364884 249372
rect 364992 249284 365172 249372
rect 365280 249284 365460 249372
rect 365714 249284 365894 249372
rect 366002 249284 366182 249372
rect 366290 249284 366470 249372
rect 366578 249284 366758 249372
rect 366866 249284 367046 249372
rect 367154 249284 367334 249372
rect 367442 249284 367622 249372
rect 367730 249284 367910 249372
rect 243214 248808 243394 248896
rect 243502 248808 243682 248896
rect 243790 248808 243970 248896
rect 244078 248808 244258 248896
rect 244366 248808 244546 248896
rect 244654 248808 244834 248896
rect 244942 248808 245122 248896
rect 245230 248808 245410 248896
rect 245664 248808 245844 248896
rect 245952 248808 246132 248896
rect 246240 248808 246420 248896
rect 246528 248808 246708 248896
rect 246816 248808 246996 248896
rect 247104 248808 247284 248896
rect 247392 248808 247572 248896
rect 247680 248808 247860 248896
rect 248114 248808 248294 248896
rect 248402 248808 248582 248896
rect 248690 248808 248870 248896
rect 248978 248808 249158 248896
rect 249266 248808 249446 248896
rect 249554 248808 249734 248896
rect 249842 248808 250022 248896
rect 250130 248808 250310 248896
rect 250564 248808 250744 248896
rect 360436 248808 360560 248896
rect 360814 248808 360994 248896
rect 361102 248808 361282 248896
rect 361390 248808 361570 248896
rect 361678 248808 361858 248896
rect 361966 248808 362146 248896
rect 362254 248808 362434 248896
rect 362542 248808 362722 248896
rect 362830 248808 363010 248896
rect 363264 248808 363444 248896
rect 363552 248808 363732 248896
rect 363840 248808 364020 248896
rect 364128 248808 364308 248896
rect 364416 248808 364596 248896
rect 364704 248808 364884 248896
rect 364992 248808 365172 248896
rect 365280 248808 365460 248896
rect 365714 248808 365894 248896
rect 366002 248808 366182 248896
rect 366290 248808 366470 248896
rect 366578 248808 366758 248896
rect 366866 248808 367046 248896
rect 367154 248808 367334 248896
rect 367442 248808 367622 248896
rect 367730 248808 367910 248896
rect 243214 248334 243394 248422
rect 243502 248334 243682 248422
rect 243790 248334 243970 248422
rect 244078 248334 244258 248422
rect 244366 248334 244546 248422
rect 244654 248334 244834 248422
rect 244942 248334 245122 248422
rect 245230 248334 245410 248422
rect 245664 248334 245844 248422
rect 245952 248334 246132 248422
rect 246240 248334 246420 248422
rect 246528 248334 246708 248422
rect 246816 248334 246996 248422
rect 247104 248334 247284 248422
rect 247392 248334 247572 248422
rect 247680 248334 247860 248422
rect 248114 248334 248294 248422
rect 248402 248334 248582 248422
rect 248690 248334 248870 248422
rect 248978 248334 249158 248422
rect 249266 248334 249446 248422
rect 249554 248334 249734 248422
rect 249842 248334 250022 248422
rect 250130 248334 250310 248422
rect 250564 248334 250744 248422
rect 360436 248334 360560 248422
rect 360814 248334 360994 248422
rect 361102 248334 361282 248422
rect 361390 248334 361570 248422
rect 361678 248334 361858 248422
rect 361966 248334 362146 248422
rect 362254 248334 362434 248422
rect 362542 248334 362722 248422
rect 362830 248334 363010 248422
rect 363264 248334 363444 248422
rect 363552 248334 363732 248422
rect 363840 248334 364020 248422
rect 364128 248334 364308 248422
rect 364416 248334 364596 248422
rect 364704 248334 364884 248422
rect 364992 248334 365172 248422
rect 365280 248334 365460 248422
rect 365714 248334 365894 248422
rect 366002 248334 366182 248422
rect 366290 248334 366470 248422
rect 366578 248334 366758 248422
rect 366866 248334 367046 248422
rect 367154 248334 367334 248422
rect 367442 248334 367622 248422
rect 367730 248334 367910 248422
rect 243214 247858 243394 247946
rect 243502 247858 243682 247946
rect 243790 247858 243970 247946
rect 244078 247858 244258 247946
rect 244366 247858 244546 247946
rect 244654 247858 244834 247946
rect 244942 247858 245122 247946
rect 245230 247858 245410 247946
rect 245664 247858 245844 247946
rect 245952 247858 246132 247946
rect 246240 247858 246420 247946
rect 246528 247858 246708 247946
rect 246816 247858 246996 247946
rect 247104 247858 247284 247946
rect 247392 247858 247572 247946
rect 247680 247858 247860 247946
rect 248114 247858 248294 247946
rect 248402 247858 248582 247946
rect 248690 247858 248870 247946
rect 248978 247858 249158 247946
rect 249266 247858 249446 247946
rect 249554 247858 249734 247946
rect 249842 247858 250022 247946
rect 250130 247858 250310 247946
rect 250564 247858 250744 247946
rect 360436 247858 360560 247946
rect 360814 247858 360994 247946
rect 361102 247858 361282 247946
rect 361390 247858 361570 247946
rect 361678 247858 361858 247946
rect 361966 247858 362146 247946
rect 362254 247858 362434 247946
rect 362542 247858 362722 247946
rect 362830 247858 363010 247946
rect 363264 247858 363444 247946
rect 363552 247858 363732 247946
rect 363840 247858 364020 247946
rect 364128 247858 364308 247946
rect 364416 247858 364596 247946
rect 364704 247858 364884 247946
rect 364992 247858 365172 247946
rect 365280 247858 365460 247946
rect 365714 247858 365894 247946
rect 366002 247858 366182 247946
rect 366290 247858 366470 247946
rect 366578 247858 366758 247946
rect 366866 247858 367046 247946
rect 367154 247858 367334 247946
rect 367442 247858 367622 247946
rect 367730 247858 367910 247946
rect 243214 247642 243394 247730
rect 243502 247642 243682 247730
rect 243790 247642 243970 247730
rect 244078 247642 244258 247730
rect 244366 247642 244546 247730
rect 244654 247642 244834 247730
rect 244942 247642 245122 247730
rect 245230 247642 245410 247730
rect 245664 247642 245844 247730
rect 245952 247642 246132 247730
rect 246240 247642 246420 247730
rect 246528 247642 246708 247730
rect 246816 247642 246996 247730
rect 247104 247642 247284 247730
rect 247392 247642 247572 247730
rect 247680 247642 247860 247730
rect 248114 247642 248294 247730
rect 248402 247642 248582 247730
rect 248690 247642 248870 247730
rect 248978 247642 249158 247730
rect 249266 247642 249446 247730
rect 249554 247642 249734 247730
rect 249842 247642 250022 247730
rect 250130 247642 250310 247730
rect 250564 247642 250744 247730
rect 360436 247642 360560 247730
rect 360814 247642 360994 247730
rect 361102 247642 361282 247730
rect 361390 247642 361570 247730
rect 361678 247642 361858 247730
rect 361966 247642 362146 247730
rect 362254 247642 362434 247730
rect 362542 247642 362722 247730
rect 362830 247642 363010 247730
rect 363264 247642 363444 247730
rect 363552 247642 363732 247730
rect 363840 247642 364020 247730
rect 364128 247642 364308 247730
rect 364416 247642 364596 247730
rect 364704 247642 364884 247730
rect 364992 247642 365172 247730
rect 365280 247642 365460 247730
rect 365714 247642 365894 247730
rect 366002 247642 366182 247730
rect 366290 247642 366470 247730
rect 366578 247642 366758 247730
rect 366866 247642 367046 247730
rect 367154 247642 367334 247730
rect 367442 247642 367622 247730
rect 367730 247642 367910 247730
rect 243214 247166 243394 247254
rect 243502 247166 243682 247254
rect 243790 247166 243970 247254
rect 244078 247166 244258 247254
rect 244366 247166 244546 247254
rect 244654 247166 244834 247254
rect 244942 247166 245122 247254
rect 245230 247166 245410 247254
rect 245664 247166 245844 247254
rect 245952 247166 246132 247254
rect 246240 247166 246420 247254
rect 246528 247166 246708 247254
rect 246816 247166 246996 247254
rect 247104 247166 247284 247254
rect 247392 247166 247572 247254
rect 247680 247166 247860 247254
rect 248114 247166 248294 247254
rect 248402 247166 248582 247254
rect 248690 247166 248870 247254
rect 248978 247166 249158 247254
rect 249266 247166 249446 247254
rect 249554 247166 249734 247254
rect 249842 247166 250022 247254
rect 250130 247166 250310 247254
rect 250564 247166 250744 247254
rect 360436 247166 360560 247254
rect 360814 247166 360994 247254
rect 361102 247166 361282 247254
rect 361390 247166 361570 247254
rect 361678 247166 361858 247254
rect 361966 247166 362146 247254
rect 362254 247166 362434 247254
rect 362542 247166 362722 247254
rect 362830 247166 363010 247254
rect 363264 247166 363444 247254
rect 363552 247166 363732 247254
rect 363840 247166 364020 247254
rect 364128 247166 364308 247254
rect 364416 247166 364596 247254
rect 364704 247166 364884 247254
rect 364992 247166 365172 247254
rect 365280 247166 365460 247254
rect 365714 247166 365894 247254
rect 366002 247166 366182 247254
rect 366290 247166 366470 247254
rect 366578 247166 366758 247254
rect 366866 247166 367046 247254
rect 367154 247166 367334 247254
rect 367442 247166 367622 247254
rect 367730 247166 367910 247254
rect 243214 246950 243394 247038
rect 243502 246950 243682 247038
rect 243790 246950 243970 247038
rect 244078 246950 244258 247038
rect 244366 246950 244546 247038
rect 244654 246950 244834 247038
rect 244942 246950 245122 247038
rect 245230 246950 245410 247038
rect 245664 246950 245844 247038
rect 245952 246950 246132 247038
rect 246240 246950 246420 247038
rect 246528 246950 246708 247038
rect 246816 246950 246996 247038
rect 247104 246950 247284 247038
rect 247392 246950 247572 247038
rect 247680 246950 247860 247038
rect 248114 246950 248294 247038
rect 248402 246950 248582 247038
rect 248690 246950 248870 247038
rect 248978 246950 249158 247038
rect 249266 246950 249446 247038
rect 249554 246950 249734 247038
rect 249842 246950 250022 247038
rect 250130 246950 250310 247038
rect 250564 246950 250744 247038
rect 360436 246950 360560 247038
rect 360814 246950 360994 247038
rect 361102 246950 361282 247038
rect 361390 246950 361570 247038
rect 361678 246950 361858 247038
rect 361966 246950 362146 247038
rect 362254 246950 362434 247038
rect 362542 246950 362722 247038
rect 362830 246950 363010 247038
rect 363264 246950 363444 247038
rect 363552 246950 363732 247038
rect 363840 246950 364020 247038
rect 364128 246950 364308 247038
rect 364416 246950 364596 247038
rect 364704 246950 364884 247038
rect 364992 246950 365172 247038
rect 365280 246950 365460 247038
rect 365714 246950 365894 247038
rect 366002 246950 366182 247038
rect 366290 246950 366470 247038
rect 366578 246950 366758 247038
rect 366866 246950 367046 247038
rect 367154 246950 367334 247038
rect 367442 246950 367622 247038
rect 367730 246950 367910 247038
rect 243214 246474 243394 246562
rect 243502 246474 243682 246562
rect 243790 246474 243970 246562
rect 244078 246474 244258 246562
rect 244366 246474 244546 246562
rect 244654 246474 244834 246562
rect 244942 246474 245122 246562
rect 245230 246474 245410 246562
rect 245664 246474 245844 246562
rect 245952 246474 246132 246562
rect 246240 246474 246420 246562
rect 246528 246474 246708 246562
rect 246816 246474 246996 246562
rect 247104 246474 247284 246562
rect 247392 246474 247572 246562
rect 247680 246474 247860 246562
rect 248114 246474 248294 246562
rect 248402 246474 248582 246562
rect 248690 246474 248870 246562
rect 248978 246474 249158 246562
rect 249266 246474 249446 246562
rect 249554 246474 249734 246562
rect 249842 246474 250022 246562
rect 250130 246474 250310 246562
rect 250564 246474 250744 246562
rect 360436 246474 360560 246562
rect 360814 246474 360994 246562
rect 361102 246474 361282 246562
rect 361390 246474 361570 246562
rect 361678 246474 361858 246562
rect 361966 246474 362146 246562
rect 362254 246474 362434 246562
rect 362542 246474 362722 246562
rect 362830 246474 363010 246562
rect 363264 246474 363444 246562
rect 363552 246474 363732 246562
rect 363840 246474 364020 246562
rect 364128 246474 364308 246562
rect 364416 246474 364596 246562
rect 364704 246474 364884 246562
rect 364992 246474 365172 246562
rect 365280 246474 365460 246562
rect 365714 246474 365894 246562
rect 366002 246474 366182 246562
rect 366290 246474 366470 246562
rect 366578 246474 366758 246562
rect 366866 246474 367046 246562
rect 367154 246474 367334 246562
rect 367442 246474 367622 246562
rect 367730 246474 367910 246562
rect 243214 246258 243394 246346
rect 243502 246258 243682 246346
rect 243790 246258 243970 246346
rect 244078 246258 244258 246346
rect 244366 246258 244546 246346
rect 244654 246258 244834 246346
rect 244942 246258 245122 246346
rect 245230 246258 245410 246346
rect 245664 246258 245844 246346
rect 245952 246258 246132 246346
rect 246240 246258 246420 246346
rect 246528 246258 246708 246346
rect 246816 246258 246996 246346
rect 247104 246258 247284 246346
rect 247392 246258 247572 246346
rect 247680 246258 247860 246346
rect 248114 246258 248294 246346
rect 248402 246258 248582 246346
rect 248690 246258 248870 246346
rect 248978 246258 249158 246346
rect 249266 246258 249446 246346
rect 249554 246258 249734 246346
rect 249842 246258 250022 246346
rect 250130 246258 250310 246346
rect 250564 246258 250744 246346
rect 360436 246258 360560 246346
rect 360814 246258 360994 246346
rect 361102 246258 361282 246346
rect 361390 246258 361570 246346
rect 361678 246258 361858 246346
rect 361966 246258 362146 246346
rect 362254 246258 362434 246346
rect 362542 246258 362722 246346
rect 362830 246258 363010 246346
rect 363264 246258 363444 246346
rect 363552 246258 363732 246346
rect 363840 246258 364020 246346
rect 364128 246258 364308 246346
rect 364416 246258 364596 246346
rect 364704 246258 364884 246346
rect 364992 246258 365172 246346
rect 365280 246258 365460 246346
rect 365714 246258 365894 246346
rect 366002 246258 366182 246346
rect 366290 246258 366470 246346
rect 366578 246258 366758 246346
rect 366866 246258 367046 246346
rect 367154 246258 367334 246346
rect 367442 246258 367622 246346
rect 367730 246258 367910 246346
rect 243214 245782 243394 245870
rect 243502 245782 243682 245870
rect 243790 245782 243970 245870
rect 244078 245782 244258 245870
rect 244366 245782 244546 245870
rect 244654 245782 244834 245870
rect 244942 245782 245122 245870
rect 245230 245782 245410 245870
rect 245664 245782 245844 245870
rect 245952 245782 246132 245870
rect 246240 245782 246420 245870
rect 246528 245782 246708 245870
rect 246816 245782 246996 245870
rect 247104 245782 247284 245870
rect 247392 245782 247572 245870
rect 247680 245782 247860 245870
rect 248114 245782 248294 245870
rect 248402 245782 248582 245870
rect 248690 245782 248870 245870
rect 248978 245782 249158 245870
rect 249266 245782 249446 245870
rect 249554 245782 249734 245870
rect 249842 245782 250022 245870
rect 250130 245782 250310 245870
rect 250564 245782 250744 245870
rect 360436 245782 360560 245870
rect 360814 245782 360994 245870
rect 361102 245782 361282 245870
rect 361390 245782 361570 245870
rect 361678 245782 361858 245870
rect 361966 245782 362146 245870
rect 362254 245782 362434 245870
rect 362542 245782 362722 245870
rect 362830 245782 363010 245870
rect 363264 245782 363444 245870
rect 363552 245782 363732 245870
rect 363840 245782 364020 245870
rect 364128 245782 364308 245870
rect 364416 245782 364596 245870
rect 364704 245782 364884 245870
rect 364992 245782 365172 245870
rect 365280 245782 365460 245870
rect 365714 245782 365894 245870
rect 366002 245782 366182 245870
rect 366290 245782 366470 245870
rect 366578 245782 366758 245870
rect 366866 245782 367046 245870
rect 367154 245782 367334 245870
rect 367442 245782 367622 245870
rect 367730 245782 367910 245870
rect 243214 245308 243394 245396
rect 243502 245308 243682 245396
rect 243790 245308 243970 245396
rect 244078 245308 244258 245396
rect 244366 245308 244546 245396
rect 244654 245308 244834 245396
rect 244942 245308 245122 245396
rect 245230 245308 245410 245396
rect 245664 245308 245844 245396
rect 245952 245308 246132 245396
rect 246240 245308 246420 245396
rect 246528 245308 246708 245396
rect 246816 245308 246996 245396
rect 247104 245308 247284 245396
rect 247392 245308 247572 245396
rect 247680 245308 247860 245396
rect 248114 245308 248294 245396
rect 248402 245308 248582 245396
rect 248690 245308 248870 245396
rect 248978 245308 249158 245396
rect 249266 245308 249446 245396
rect 249554 245308 249734 245396
rect 249842 245308 250022 245396
rect 250130 245308 250310 245396
rect 250564 245308 250744 245396
rect 360436 245308 360560 245396
rect 360814 245308 360994 245396
rect 361102 245308 361282 245396
rect 361390 245308 361570 245396
rect 361678 245308 361858 245396
rect 361966 245308 362146 245396
rect 362254 245308 362434 245396
rect 362542 245308 362722 245396
rect 362830 245308 363010 245396
rect 363264 245308 363444 245396
rect 363552 245308 363732 245396
rect 363840 245308 364020 245396
rect 364128 245308 364308 245396
rect 364416 245308 364596 245396
rect 364704 245308 364884 245396
rect 364992 245308 365172 245396
rect 365280 245308 365460 245396
rect 365714 245308 365894 245396
rect 366002 245308 366182 245396
rect 366290 245308 366470 245396
rect 366578 245308 366758 245396
rect 366866 245308 367046 245396
rect 367154 245308 367334 245396
rect 367442 245308 367622 245396
rect 367730 245308 367910 245396
rect 243214 244832 243394 244920
rect 243502 244832 243682 244920
rect 243790 244832 243970 244920
rect 244078 244832 244258 244920
rect 244366 244832 244546 244920
rect 244654 244832 244834 244920
rect 244942 244832 245122 244920
rect 245230 244832 245410 244920
rect 245664 244832 245844 244920
rect 245952 244832 246132 244920
rect 246240 244832 246420 244920
rect 246528 244832 246708 244920
rect 246816 244832 246996 244920
rect 247104 244832 247284 244920
rect 247392 244832 247572 244920
rect 247680 244832 247860 244920
rect 248114 244832 248294 244920
rect 248402 244832 248582 244920
rect 248690 244832 248870 244920
rect 248978 244832 249158 244920
rect 249266 244832 249446 244920
rect 249554 244832 249734 244920
rect 249842 244832 250022 244920
rect 250130 244832 250310 244920
rect 250564 244832 250744 244920
rect 360436 244832 360560 244920
rect 360814 244832 360994 244920
rect 361102 244832 361282 244920
rect 361390 244832 361570 244920
rect 361678 244832 361858 244920
rect 361966 244832 362146 244920
rect 362254 244832 362434 244920
rect 362542 244832 362722 244920
rect 362830 244832 363010 244920
rect 363264 244832 363444 244920
rect 363552 244832 363732 244920
rect 363840 244832 364020 244920
rect 364128 244832 364308 244920
rect 364416 244832 364596 244920
rect 364704 244832 364884 244920
rect 364992 244832 365172 244920
rect 365280 244832 365460 244920
rect 365714 244832 365894 244920
rect 366002 244832 366182 244920
rect 366290 244832 366470 244920
rect 366578 244832 366758 244920
rect 366866 244832 367046 244920
rect 367154 244832 367334 244920
rect 367442 244832 367622 244920
rect 367730 244832 367910 244920
rect 243214 244616 243394 244704
rect 243502 244616 243682 244704
rect 243790 244616 243970 244704
rect 244078 244616 244258 244704
rect 244366 244616 244546 244704
rect 244654 244616 244834 244704
rect 244942 244616 245122 244704
rect 245230 244616 245410 244704
rect 245664 244616 245844 244704
rect 245952 244616 246132 244704
rect 246240 244616 246420 244704
rect 246528 244616 246708 244704
rect 246816 244616 246996 244704
rect 247104 244616 247284 244704
rect 247392 244616 247572 244704
rect 247680 244616 247860 244704
rect 248114 244616 248294 244704
rect 248402 244616 248582 244704
rect 248690 244616 248870 244704
rect 248978 244616 249158 244704
rect 249266 244616 249446 244704
rect 249554 244616 249734 244704
rect 249842 244616 250022 244704
rect 250130 244616 250310 244704
rect 250564 244616 250744 244704
rect 360436 244616 360560 244704
rect 360814 244616 360994 244704
rect 361102 244616 361282 244704
rect 361390 244616 361570 244704
rect 361678 244616 361858 244704
rect 361966 244616 362146 244704
rect 362254 244616 362434 244704
rect 362542 244616 362722 244704
rect 362830 244616 363010 244704
rect 363264 244616 363444 244704
rect 363552 244616 363732 244704
rect 363840 244616 364020 244704
rect 364128 244616 364308 244704
rect 364416 244616 364596 244704
rect 364704 244616 364884 244704
rect 364992 244616 365172 244704
rect 365280 244616 365460 244704
rect 365714 244616 365894 244704
rect 366002 244616 366182 244704
rect 366290 244616 366470 244704
rect 366578 244616 366758 244704
rect 366866 244616 367046 244704
rect 367154 244616 367334 244704
rect 367442 244616 367622 244704
rect 367730 244616 367910 244704
rect 243214 244140 243394 244228
rect 243502 244140 243682 244228
rect 243790 244140 243970 244228
rect 244078 244140 244258 244228
rect 244366 244140 244546 244228
rect 244654 244140 244834 244228
rect 244942 244140 245122 244228
rect 245230 244140 245410 244228
rect 245664 244140 245844 244228
rect 245952 244140 246132 244228
rect 246240 244140 246420 244228
rect 246528 244140 246708 244228
rect 246816 244140 246996 244228
rect 247104 244140 247284 244228
rect 247392 244140 247572 244228
rect 247680 244140 247860 244228
rect 248114 244140 248294 244228
rect 248402 244140 248582 244228
rect 248690 244140 248870 244228
rect 248978 244140 249158 244228
rect 249266 244140 249446 244228
rect 249554 244140 249734 244228
rect 249842 244140 250022 244228
rect 250130 244140 250310 244228
rect 250564 244140 250744 244228
rect 360436 244140 360560 244228
rect 360814 244140 360994 244228
rect 361102 244140 361282 244228
rect 361390 244140 361570 244228
rect 361678 244140 361858 244228
rect 361966 244140 362146 244228
rect 362254 244140 362434 244228
rect 362542 244140 362722 244228
rect 362830 244140 363010 244228
rect 363264 244140 363444 244228
rect 363552 244140 363732 244228
rect 363840 244140 364020 244228
rect 364128 244140 364308 244228
rect 364416 244140 364596 244228
rect 364704 244140 364884 244228
rect 364992 244140 365172 244228
rect 365280 244140 365460 244228
rect 365714 244140 365894 244228
rect 366002 244140 366182 244228
rect 366290 244140 366470 244228
rect 366578 244140 366758 244228
rect 366866 244140 367046 244228
rect 367154 244140 367334 244228
rect 367442 244140 367622 244228
rect 367730 244140 367910 244228
rect 243214 243924 243394 244012
rect 243502 243924 243682 244012
rect 243790 243924 243970 244012
rect 244078 243924 244258 244012
rect 244366 243924 244546 244012
rect 244654 243924 244834 244012
rect 244942 243924 245122 244012
rect 245230 243924 245410 244012
rect 245664 243924 245844 244012
rect 245952 243924 246132 244012
rect 246240 243924 246420 244012
rect 246528 243924 246708 244012
rect 246816 243924 246996 244012
rect 247104 243924 247284 244012
rect 247392 243924 247572 244012
rect 247680 243924 247860 244012
rect 248114 243924 248294 244012
rect 248402 243924 248582 244012
rect 248690 243924 248870 244012
rect 248978 243924 249158 244012
rect 249266 243924 249446 244012
rect 249554 243924 249734 244012
rect 249842 243924 250022 244012
rect 250130 243924 250310 244012
rect 250564 243924 250744 244012
rect 360436 243924 360560 244012
rect 360814 243924 360994 244012
rect 361102 243924 361282 244012
rect 361390 243924 361570 244012
rect 361678 243924 361858 244012
rect 361966 243924 362146 244012
rect 362254 243924 362434 244012
rect 362542 243924 362722 244012
rect 362830 243924 363010 244012
rect 363264 243924 363444 244012
rect 363552 243924 363732 244012
rect 363840 243924 364020 244012
rect 364128 243924 364308 244012
rect 364416 243924 364596 244012
rect 364704 243924 364884 244012
rect 364992 243924 365172 244012
rect 365280 243924 365460 244012
rect 365714 243924 365894 244012
rect 366002 243924 366182 244012
rect 366290 243924 366470 244012
rect 366578 243924 366758 244012
rect 366866 243924 367046 244012
rect 367154 243924 367334 244012
rect 367442 243924 367622 244012
rect 367730 243924 367910 244012
rect 243214 243448 243394 243536
rect 243502 243448 243682 243536
rect 243790 243448 243970 243536
rect 244078 243448 244258 243536
rect 244366 243448 244546 243536
rect 244654 243448 244834 243536
rect 244942 243448 245122 243536
rect 245230 243448 245410 243536
rect 245664 243448 245844 243536
rect 245952 243448 246132 243536
rect 246240 243448 246420 243536
rect 246528 243448 246708 243536
rect 246816 243448 246996 243536
rect 247104 243448 247284 243536
rect 247392 243448 247572 243536
rect 247680 243448 247860 243536
rect 248114 243448 248294 243536
rect 248402 243448 248582 243536
rect 248690 243448 248870 243536
rect 248978 243448 249158 243536
rect 249266 243448 249446 243536
rect 249554 243448 249734 243536
rect 249842 243448 250022 243536
rect 250130 243448 250310 243536
rect 250564 243448 250744 243536
rect 360436 243448 360560 243536
rect 360814 243448 360994 243536
rect 361102 243448 361282 243536
rect 361390 243448 361570 243536
rect 361678 243448 361858 243536
rect 361966 243448 362146 243536
rect 362254 243448 362434 243536
rect 362542 243448 362722 243536
rect 362830 243448 363010 243536
rect 363264 243448 363444 243536
rect 363552 243448 363732 243536
rect 363840 243448 364020 243536
rect 364128 243448 364308 243536
rect 364416 243448 364596 243536
rect 364704 243448 364884 243536
rect 364992 243448 365172 243536
rect 365280 243448 365460 243536
rect 365714 243448 365894 243536
rect 366002 243448 366182 243536
rect 366290 243448 366470 243536
rect 366578 243448 366758 243536
rect 366866 243448 367046 243536
rect 367154 243448 367334 243536
rect 367442 243448 367622 243536
rect 367730 243448 367910 243536
rect 243214 243232 243394 243320
rect 243502 243232 243682 243320
rect 243790 243232 243970 243320
rect 244078 243232 244258 243320
rect 244366 243232 244546 243320
rect 244654 243232 244834 243320
rect 244942 243232 245122 243320
rect 245230 243232 245410 243320
rect 245664 243232 245844 243320
rect 245952 243232 246132 243320
rect 246240 243232 246420 243320
rect 246528 243232 246708 243320
rect 246816 243232 246996 243320
rect 247104 243232 247284 243320
rect 247392 243232 247572 243320
rect 247680 243232 247860 243320
rect 248114 243232 248294 243320
rect 248402 243232 248582 243320
rect 248690 243232 248870 243320
rect 248978 243232 249158 243320
rect 249266 243232 249446 243320
rect 249554 243232 249734 243320
rect 249842 243232 250022 243320
rect 250130 243232 250310 243320
rect 250564 243232 250744 243320
rect 360436 243232 360560 243320
rect 360814 243232 360994 243320
rect 361102 243232 361282 243320
rect 361390 243232 361570 243320
rect 361678 243232 361858 243320
rect 361966 243232 362146 243320
rect 362254 243232 362434 243320
rect 362542 243232 362722 243320
rect 362830 243232 363010 243320
rect 363264 243232 363444 243320
rect 363552 243232 363732 243320
rect 363840 243232 364020 243320
rect 364128 243232 364308 243320
rect 364416 243232 364596 243320
rect 364704 243232 364884 243320
rect 364992 243232 365172 243320
rect 365280 243232 365460 243320
rect 365714 243232 365894 243320
rect 366002 243232 366182 243320
rect 366290 243232 366470 243320
rect 366578 243232 366758 243320
rect 366866 243232 367046 243320
rect 367154 243232 367334 243320
rect 367442 243232 367622 243320
rect 367730 243232 367910 243320
rect 243214 242756 243394 242844
rect 243502 242756 243682 242844
rect 243790 242756 243970 242844
rect 244078 242756 244258 242844
rect 244366 242756 244546 242844
rect 244654 242756 244834 242844
rect 244942 242756 245122 242844
rect 245230 242756 245410 242844
rect 245664 242756 245844 242844
rect 245952 242756 246132 242844
rect 246240 242756 246420 242844
rect 246528 242756 246708 242844
rect 246816 242756 246996 242844
rect 247104 242756 247284 242844
rect 247392 242756 247572 242844
rect 247680 242756 247860 242844
rect 248114 242756 248294 242844
rect 248402 242756 248582 242844
rect 248690 242756 248870 242844
rect 248978 242756 249158 242844
rect 249266 242756 249446 242844
rect 249554 242756 249734 242844
rect 249842 242756 250022 242844
rect 250130 242756 250310 242844
rect 250564 242756 250744 242844
rect 360436 242756 360560 242844
rect 360814 242756 360994 242844
rect 361102 242756 361282 242844
rect 361390 242756 361570 242844
rect 361678 242756 361858 242844
rect 361966 242756 362146 242844
rect 362254 242756 362434 242844
rect 362542 242756 362722 242844
rect 362830 242756 363010 242844
rect 363264 242756 363444 242844
rect 363552 242756 363732 242844
rect 363840 242756 364020 242844
rect 364128 242756 364308 242844
rect 364416 242756 364596 242844
rect 364704 242756 364884 242844
rect 364992 242756 365172 242844
rect 365280 242756 365460 242844
rect 365714 242756 365894 242844
rect 366002 242756 366182 242844
rect 366290 242756 366470 242844
rect 366578 242756 366758 242844
rect 366866 242756 367046 242844
rect 367154 242756 367334 242844
rect 367442 242756 367622 242844
rect 367730 242756 367910 242844
rect 243214 242282 243394 242370
rect 243502 242282 243682 242370
rect 243790 242282 243970 242370
rect 244078 242282 244258 242370
rect 244366 242282 244546 242370
rect 244654 242282 244834 242370
rect 244942 242282 245122 242370
rect 245230 242282 245410 242370
rect 245664 242282 245844 242370
rect 245952 242282 246132 242370
rect 246240 242282 246420 242370
rect 246528 242282 246708 242370
rect 246816 242282 246996 242370
rect 247104 242282 247284 242370
rect 247392 242282 247572 242370
rect 247680 242282 247860 242370
rect 248114 242282 248294 242370
rect 248402 242282 248582 242370
rect 248690 242282 248870 242370
rect 248978 242282 249158 242370
rect 249266 242282 249446 242370
rect 249554 242282 249734 242370
rect 249842 242282 250022 242370
rect 250130 242282 250310 242370
rect 250564 242282 250744 242370
rect 360436 242282 360560 242370
rect 360814 242282 360994 242370
rect 361102 242282 361282 242370
rect 361390 242282 361570 242370
rect 361678 242282 361858 242370
rect 361966 242282 362146 242370
rect 362254 242282 362434 242370
rect 362542 242282 362722 242370
rect 362830 242282 363010 242370
rect 363264 242282 363444 242370
rect 363552 242282 363732 242370
rect 363840 242282 364020 242370
rect 364128 242282 364308 242370
rect 364416 242282 364596 242370
rect 364704 242282 364884 242370
rect 364992 242282 365172 242370
rect 365280 242282 365460 242370
rect 365714 242282 365894 242370
rect 366002 242282 366182 242370
rect 366290 242282 366470 242370
rect 366578 242282 366758 242370
rect 366866 242282 367046 242370
rect 367154 242282 367334 242370
rect 367442 242282 367622 242370
rect 367730 242282 367910 242370
rect 243214 241806 243394 241894
rect 243502 241806 243682 241894
rect 243790 241806 243970 241894
rect 244078 241806 244258 241894
rect 244366 241806 244546 241894
rect 244654 241806 244834 241894
rect 244942 241806 245122 241894
rect 245230 241806 245410 241894
rect 245664 241806 245844 241894
rect 245952 241806 246132 241894
rect 246240 241806 246420 241894
rect 246528 241806 246708 241894
rect 246816 241806 246996 241894
rect 247104 241806 247284 241894
rect 247392 241806 247572 241894
rect 247680 241806 247860 241894
rect 248114 241806 248294 241894
rect 248402 241806 248582 241894
rect 248690 241806 248870 241894
rect 248978 241806 249158 241894
rect 249266 241806 249446 241894
rect 249554 241806 249734 241894
rect 249842 241806 250022 241894
rect 250130 241806 250310 241894
rect 250564 241806 250744 241894
rect 360436 241806 360560 241894
rect 360814 241806 360994 241894
rect 361102 241806 361282 241894
rect 361390 241806 361570 241894
rect 361678 241806 361858 241894
rect 361966 241806 362146 241894
rect 362254 241806 362434 241894
rect 362542 241806 362722 241894
rect 362830 241806 363010 241894
rect 363264 241806 363444 241894
rect 363552 241806 363732 241894
rect 363840 241806 364020 241894
rect 364128 241806 364308 241894
rect 364416 241806 364596 241894
rect 364704 241806 364884 241894
rect 364992 241806 365172 241894
rect 365280 241806 365460 241894
rect 365714 241806 365894 241894
rect 366002 241806 366182 241894
rect 366290 241806 366470 241894
rect 366578 241806 366758 241894
rect 366866 241806 367046 241894
rect 367154 241806 367334 241894
rect 367442 241806 367622 241894
rect 367730 241806 367910 241894
rect 243214 241590 243394 241678
rect 243502 241590 243682 241678
rect 243790 241590 243970 241678
rect 244078 241590 244258 241678
rect 244366 241590 244546 241678
rect 244654 241590 244834 241678
rect 244942 241590 245122 241678
rect 245230 241590 245410 241678
rect 245664 241590 245844 241678
rect 245952 241590 246132 241678
rect 246240 241590 246420 241678
rect 246528 241590 246708 241678
rect 246816 241590 246996 241678
rect 247104 241590 247284 241678
rect 247392 241590 247572 241678
rect 247680 241590 247860 241678
rect 248114 241590 248294 241678
rect 248402 241590 248582 241678
rect 248690 241590 248870 241678
rect 248978 241590 249158 241678
rect 249266 241590 249446 241678
rect 249554 241590 249734 241678
rect 249842 241590 250022 241678
rect 250130 241590 250310 241678
rect 250564 241590 250744 241678
rect 360436 241590 360560 241678
rect 360814 241590 360994 241678
rect 361102 241590 361282 241678
rect 361390 241590 361570 241678
rect 361678 241590 361858 241678
rect 361966 241590 362146 241678
rect 362254 241590 362434 241678
rect 362542 241590 362722 241678
rect 362830 241590 363010 241678
rect 363264 241590 363444 241678
rect 363552 241590 363732 241678
rect 363840 241590 364020 241678
rect 364128 241590 364308 241678
rect 364416 241590 364596 241678
rect 364704 241590 364884 241678
rect 364992 241590 365172 241678
rect 365280 241590 365460 241678
rect 365714 241590 365894 241678
rect 366002 241590 366182 241678
rect 366290 241590 366470 241678
rect 366578 241590 366758 241678
rect 366866 241590 367046 241678
rect 367154 241590 367334 241678
rect 367442 241590 367622 241678
rect 367730 241590 367910 241678
rect 243214 241114 243394 241202
rect 243502 241114 243682 241202
rect 243790 241114 243970 241202
rect 244078 241114 244258 241202
rect 244366 241114 244546 241202
rect 244654 241114 244834 241202
rect 244942 241114 245122 241202
rect 245230 241114 245410 241202
rect 245664 241114 245844 241202
rect 245952 241114 246132 241202
rect 246240 241114 246420 241202
rect 246528 241114 246708 241202
rect 246816 241114 246996 241202
rect 247104 241114 247284 241202
rect 247392 241114 247572 241202
rect 247680 241114 247860 241202
rect 248114 241114 248294 241202
rect 248402 241114 248582 241202
rect 248690 241114 248870 241202
rect 248978 241114 249158 241202
rect 249266 241114 249446 241202
rect 249554 241114 249734 241202
rect 249842 241114 250022 241202
rect 250130 241114 250310 241202
rect 250564 241114 250744 241202
rect 360436 241114 360560 241202
rect 360814 241114 360994 241202
rect 361102 241114 361282 241202
rect 361390 241114 361570 241202
rect 361678 241114 361858 241202
rect 361966 241114 362146 241202
rect 362254 241114 362434 241202
rect 362542 241114 362722 241202
rect 362830 241114 363010 241202
rect 363264 241114 363444 241202
rect 363552 241114 363732 241202
rect 363840 241114 364020 241202
rect 364128 241114 364308 241202
rect 364416 241114 364596 241202
rect 364704 241114 364884 241202
rect 364992 241114 365172 241202
rect 365280 241114 365460 241202
rect 365714 241114 365894 241202
rect 366002 241114 366182 241202
rect 366290 241114 366470 241202
rect 366578 241114 366758 241202
rect 366866 241114 367046 241202
rect 367154 241114 367334 241202
rect 367442 241114 367622 241202
rect 367730 241114 367910 241202
rect 243214 240898 243394 240986
rect 243502 240898 243682 240986
rect 243790 240898 243970 240986
rect 244078 240898 244258 240986
rect 244366 240898 244546 240986
rect 244654 240898 244834 240986
rect 244942 240898 245122 240986
rect 245230 240898 245410 240986
rect 245664 240898 245844 240986
rect 245952 240898 246132 240986
rect 246240 240898 246420 240986
rect 246528 240898 246708 240986
rect 246816 240898 246996 240986
rect 247104 240898 247284 240986
rect 247392 240898 247572 240986
rect 247680 240898 247860 240986
rect 248114 240898 248294 240986
rect 248402 240898 248582 240986
rect 248690 240898 248870 240986
rect 248978 240898 249158 240986
rect 249266 240898 249446 240986
rect 249554 240898 249734 240986
rect 249842 240898 250022 240986
rect 250130 240898 250310 240986
rect 250564 240898 250744 240986
rect 360436 240898 360560 240986
rect 360814 240898 360994 240986
rect 361102 240898 361282 240986
rect 361390 240898 361570 240986
rect 361678 240898 361858 240986
rect 361966 240898 362146 240986
rect 362254 240898 362434 240986
rect 362542 240898 362722 240986
rect 362830 240898 363010 240986
rect 363264 240898 363444 240986
rect 363552 240898 363732 240986
rect 363840 240898 364020 240986
rect 364128 240898 364308 240986
rect 364416 240898 364596 240986
rect 364704 240898 364884 240986
rect 364992 240898 365172 240986
rect 365280 240898 365460 240986
rect 365714 240898 365894 240986
rect 366002 240898 366182 240986
rect 366290 240898 366470 240986
rect 366578 240898 366758 240986
rect 366866 240898 367046 240986
rect 367154 240898 367334 240986
rect 367442 240898 367622 240986
rect 367730 240898 367910 240986
rect 243214 240422 243394 240510
rect 243502 240422 243682 240510
rect 243790 240422 243970 240510
rect 244078 240422 244258 240510
rect 244366 240422 244546 240510
rect 244654 240422 244834 240510
rect 244942 240422 245122 240510
rect 245230 240422 245410 240510
rect 245664 240422 245844 240510
rect 245952 240422 246132 240510
rect 246240 240422 246420 240510
rect 246528 240422 246708 240510
rect 246816 240422 246996 240510
rect 247104 240422 247284 240510
rect 247392 240422 247572 240510
rect 247680 240422 247860 240510
rect 248114 240422 248294 240510
rect 248402 240422 248582 240510
rect 248690 240422 248870 240510
rect 248978 240422 249158 240510
rect 249266 240422 249446 240510
rect 249554 240422 249734 240510
rect 249842 240422 250022 240510
rect 250130 240422 250310 240510
rect 250564 240422 250744 240510
rect 360436 240422 360560 240510
rect 360814 240422 360994 240510
rect 361102 240422 361282 240510
rect 361390 240422 361570 240510
rect 361678 240422 361858 240510
rect 361966 240422 362146 240510
rect 362254 240422 362434 240510
rect 362542 240422 362722 240510
rect 362830 240422 363010 240510
rect 363264 240422 363444 240510
rect 363552 240422 363732 240510
rect 363840 240422 364020 240510
rect 364128 240422 364308 240510
rect 364416 240422 364596 240510
rect 364704 240422 364884 240510
rect 364992 240422 365172 240510
rect 365280 240422 365460 240510
rect 365714 240422 365894 240510
rect 366002 240422 366182 240510
rect 366290 240422 366470 240510
rect 366578 240422 366758 240510
rect 366866 240422 367046 240510
rect 367154 240422 367334 240510
rect 367442 240422 367622 240510
rect 367730 240422 367910 240510
rect 243214 240206 243394 240294
rect 243502 240206 243682 240294
rect 243790 240206 243970 240294
rect 244078 240206 244258 240294
rect 244366 240206 244546 240294
rect 244654 240206 244834 240294
rect 244942 240206 245122 240294
rect 245230 240206 245410 240294
rect 245664 240206 245844 240294
rect 245952 240206 246132 240294
rect 246240 240206 246420 240294
rect 246528 240206 246708 240294
rect 246816 240206 246996 240294
rect 247104 240206 247284 240294
rect 247392 240206 247572 240294
rect 247680 240206 247860 240294
rect 248114 240206 248294 240294
rect 248402 240206 248582 240294
rect 248690 240206 248870 240294
rect 248978 240206 249158 240294
rect 249266 240206 249446 240294
rect 249554 240206 249734 240294
rect 249842 240206 250022 240294
rect 250130 240206 250310 240294
rect 250564 240206 250744 240294
rect 360436 240206 360560 240294
rect 360814 240206 360994 240294
rect 361102 240206 361282 240294
rect 361390 240206 361570 240294
rect 361678 240206 361858 240294
rect 361966 240206 362146 240294
rect 362254 240206 362434 240294
rect 362542 240206 362722 240294
rect 362830 240206 363010 240294
rect 363264 240206 363444 240294
rect 363552 240206 363732 240294
rect 363840 240206 364020 240294
rect 364128 240206 364308 240294
rect 364416 240206 364596 240294
rect 364704 240206 364884 240294
rect 364992 240206 365172 240294
rect 365280 240206 365460 240294
rect 365714 240206 365894 240294
rect 366002 240206 366182 240294
rect 366290 240206 366470 240294
rect 366578 240206 366758 240294
rect 366866 240206 367046 240294
rect 367154 240206 367334 240294
rect 367442 240206 367622 240294
rect 367730 240206 367910 240294
rect 243214 239730 243394 239818
rect 243502 239730 243682 239818
rect 243790 239730 243970 239818
rect 244078 239730 244258 239818
rect 244366 239730 244546 239818
rect 244654 239730 244834 239818
rect 244942 239730 245122 239818
rect 245230 239730 245410 239818
rect 245664 239730 245844 239818
rect 245952 239730 246132 239818
rect 246240 239730 246420 239818
rect 246528 239730 246708 239818
rect 246816 239730 246996 239818
rect 247104 239730 247284 239818
rect 247392 239730 247572 239818
rect 247680 239730 247860 239818
rect 248114 239730 248294 239818
rect 248402 239730 248582 239818
rect 248690 239730 248870 239818
rect 248978 239730 249158 239818
rect 249266 239730 249446 239818
rect 249554 239730 249734 239818
rect 249842 239730 250022 239818
rect 250130 239730 250310 239818
rect 250564 239730 250744 239818
rect 360436 239730 360560 239818
rect 360814 239730 360994 239818
rect 361102 239730 361282 239818
rect 361390 239730 361570 239818
rect 361678 239730 361858 239818
rect 361966 239730 362146 239818
rect 362254 239730 362434 239818
rect 362542 239730 362722 239818
rect 362830 239730 363010 239818
rect 363264 239730 363444 239818
rect 363552 239730 363732 239818
rect 363840 239730 364020 239818
rect 364128 239730 364308 239818
rect 364416 239730 364596 239818
rect 364704 239730 364884 239818
rect 364992 239730 365172 239818
rect 365280 239730 365460 239818
rect 365714 239730 365894 239818
rect 366002 239730 366182 239818
rect 366290 239730 366470 239818
rect 366578 239730 366758 239818
rect 366866 239730 367046 239818
rect 367154 239730 367334 239818
rect 367442 239730 367622 239818
rect 367730 239730 367910 239818
rect 243214 239256 243394 239344
rect 243502 239256 243682 239344
rect 243790 239256 243970 239344
rect 244078 239256 244258 239344
rect 244366 239256 244546 239344
rect 244654 239256 244834 239344
rect 244942 239256 245122 239344
rect 245230 239256 245410 239344
rect 245664 239256 245844 239344
rect 245952 239256 246132 239344
rect 246240 239256 246420 239344
rect 246528 239256 246708 239344
rect 246816 239256 246996 239344
rect 247104 239256 247284 239344
rect 247392 239256 247572 239344
rect 247680 239256 247860 239344
rect 248114 239256 248294 239344
rect 248402 239256 248582 239344
rect 248690 239256 248870 239344
rect 248978 239256 249158 239344
rect 249266 239256 249446 239344
rect 249554 239256 249734 239344
rect 249842 239256 250022 239344
rect 250130 239256 250310 239344
rect 250564 239256 250744 239344
rect 360436 239256 360560 239344
rect 360814 239256 360994 239344
rect 361102 239256 361282 239344
rect 361390 239256 361570 239344
rect 361678 239256 361858 239344
rect 361966 239256 362146 239344
rect 362254 239256 362434 239344
rect 362542 239256 362722 239344
rect 362830 239256 363010 239344
rect 363264 239256 363444 239344
rect 363552 239256 363732 239344
rect 363840 239256 364020 239344
rect 364128 239256 364308 239344
rect 364416 239256 364596 239344
rect 364704 239256 364884 239344
rect 364992 239256 365172 239344
rect 365280 239256 365460 239344
rect 365714 239256 365894 239344
rect 366002 239256 366182 239344
rect 366290 239256 366470 239344
rect 366578 239256 366758 239344
rect 366866 239256 367046 239344
rect 367154 239256 367334 239344
rect 367442 239256 367622 239344
rect 367730 239256 367910 239344
rect 243214 238780 243394 238868
rect 243502 238780 243682 238868
rect 243790 238780 243970 238868
rect 244078 238780 244258 238868
rect 244366 238780 244546 238868
rect 244654 238780 244834 238868
rect 244942 238780 245122 238868
rect 245230 238780 245410 238868
rect 245664 238780 245844 238868
rect 245952 238780 246132 238868
rect 246240 238780 246420 238868
rect 246528 238780 246708 238868
rect 246816 238780 246996 238868
rect 247104 238780 247284 238868
rect 247392 238780 247572 238868
rect 247680 238780 247860 238868
rect 248114 238780 248294 238868
rect 248402 238780 248582 238868
rect 248690 238780 248870 238868
rect 248978 238780 249158 238868
rect 249266 238780 249446 238868
rect 249554 238780 249734 238868
rect 249842 238780 250022 238868
rect 250130 238780 250310 238868
rect 250564 238780 250744 238868
rect 360436 238780 360560 238868
rect 360814 238780 360994 238868
rect 361102 238780 361282 238868
rect 361390 238780 361570 238868
rect 361678 238780 361858 238868
rect 361966 238780 362146 238868
rect 362254 238780 362434 238868
rect 362542 238780 362722 238868
rect 362830 238780 363010 238868
rect 363264 238780 363444 238868
rect 363552 238780 363732 238868
rect 363840 238780 364020 238868
rect 364128 238780 364308 238868
rect 364416 238780 364596 238868
rect 364704 238780 364884 238868
rect 364992 238780 365172 238868
rect 365280 238780 365460 238868
rect 365714 238780 365894 238868
rect 366002 238780 366182 238868
rect 366290 238780 366470 238868
rect 366578 238780 366758 238868
rect 366866 238780 367046 238868
rect 367154 238780 367334 238868
rect 367442 238780 367622 238868
rect 367730 238780 367910 238868
rect 243214 238564 243394 238652
rect 243502 238564 243682 238652
rect 243790 238564 243970 238652
rect 244078 238564 244258 238652
rect 244366 238564 244546 238652
rect 244654 238564 244834 238652
rect 244942 238564 245122 238652
rect 245230 238564 245410 238652
rect 245664 238564 245844 238652
rect 245952 238564 246132 238652
rect 246240 238564 246420 238652
rect 246528 238564 246708 238652
rect 246816 238564 246996 238652
rect 247104 238564 247284 238652
rect 247392 238564 247572 238652
rect 247680 238564 247860 238652
rect 248114 238564 248294 238652
rect 248402 238564 248582 238652
rect 248690 238564 248870 238652
rect 248978 238564 249158 238652
rect 249266 238564 249446 238652
rect 249554 238564 249734 238652
rect 249842 238564 250022 238652
rect 250130 238564 250310 238652
rect 250564 238564 250744 238652
rect 360436 238564 360560 238652
rect 360814 238564 360994 238652
rect 361102 238564 361282 238652
rect 361390 238564 361570 238652
rect 361678 238564 361858 238652
rect 361966 238564 362146 238652
rect 362254 238564 362434 238652
rect 362542 238564 362722 238652
rect 362830 238564 363010 238652
rect 363264 238564 363444 238652
rect 363552 238564 363732 238652
rect 363840 238564 364020 238652
rect 364128 238564 364308 238652
rect 364416 238564 364596 238652
rect 364704 238564 364884 238652
rect 364992 238564 365172 238652
rect 365280 238564 365460 238652
rect 365714 238564 365894 238652
rect 366002 238564 366182 238652
rect 366290 238564 366470 238652
rect 366578 238564 366758 238652
rect 366866 238564 367046 238652
rect 367154 238564 367334 238652
rect 367442 238564 367622 238652
rect 367730 238564 367910 238652
rect 243214 238088 243394 238176
rect 243502 238088 243682 238176
rect 243790 238088 243970 238176
rect 244078 238088 244258 238176
rect 244366 238088 244546 238176
rect 244654 238088 244834 238176
rect 244942 238088 245122 238176
rect 245230 238088 245410 238176
rect 245664 238088 245844 238176
rect 245952 238088 246132 238176
rect 246240 238088 246420 238176
rect 246528 238088 246708 238176
rect 246816 238088 246996 238176
rect 247104 238088 247284 238176
rect 247392 238088 247572 238176
rect 247680 238088 247860 238176
rect 248114 238088 248294 238176
rect 248402 238088 248582 238176
rect 248690 238088 248870 238176
rect 248978 238088 249158 238176
rect 249266 238088 249446 238176
rect 249554 238088 249734 238176
rect 249842 238088 250022 238176
rect 250130 238088 250310 238176
rect 250564 238088 250744 238176
rect 360436 238088 360560 238176
rect 360814 238088 360994 238176
rect 361102 238088 361282 238176
rect 361390 238088 361570 238176
rect 361678 238088 361858 238176
rect 361966 238088 362146 238176
rect 362254 238088 362434 238176
rect 362542 238088 362722 238176
rect 362830 238088 363010 238176
rect 363264 238088 363444 238176
rect 363552 238088 363732 238176
rect 363840 238088 364020 238176
rect 364128 238088 364308 238176
rect 364416 238088 364596 238176
rect 364704 238088 364884 238176
rect 364992 238088 365172 238176
rect 365280 238088 365460 238176
rect 365714 238088 365894 238176
rect 366002 238088 366182 238176
rect 366290 238088 366470 238176
rect 366578 238088 366758 238176
rect 366866 238088 367046 238176
rect 367154 238088 367334 238176
rect 367442 238088 367622 238176
rect 367730 238088 367910 238176
rect 243214 237872 243394 237960
rect 243502 237872 243682 237960
rect 243790 237872 243970 237960
rect 244078 237872 244258 237960
rect 244366 237872 244546 237960
rect 244654 237872 244834 237960
rect 244942 237872 245122 237960
rect 245230 237872 245410 237960
rect 245664 237872 245844 237960
rect 245952 237872 246132 237960
rect 246240 237872 246420 237960
rect 246528 237872 246708 237960
rect 246816 237872 246996 237960
rect 247104 237872 247284 237960
rect 247392 237872 247572 237960
rect 247680 237872 247860 237960
rect 248114 237872 248294 237960
rect 248402 237872 248582 237960
rect 248690 237872 248870 237960
rect 248978 237872 249158 237960
rect 249266 237872 249446 237960
rect 249554 237872 249734 237960
rect 249842 237872 250022 237960
rect 250130 237872 250310 237960
rect 250564 237872 250744 237960
rect 360436 237872 360560 237960
rect 360814 237872 360994 237960
rect 361102 237872 361282 237960
rect 361390 237872 361570 237960
rect 361678 237872 361858 237960
rect 361966 237872 362146 237960
rect 362254 237872 362434 237960
rect 362542 237872 362722 237960
rect 362830 237872 363010 237960
rect 363264 237872 363444 237960
rect 363552 237872 363732 237960
rect 363840 237872 364020 237960
rect 364128 237872 364308 237960
rect 364416 237872 364596 237960
rect 364704 237872 364884 237960
rect 364992 237872 365172 237960
rect 365280 237872 365460 237960
rect 365714 237872 365894 237960
rect 366002 237872 366182 237960
rect 366290 237872 366470 237960
rect 366578 237872 366758 237960
rect 366866 237872 367046 237960
rect 367154 237872 367334 237960
rect 367442 237872 367622 237960
rect 367730 237872 367910 237960
rect 243214 237396 243394 237484
rect 243502 237396 243682 237484
rect 243790 237396 243970 237484
rect 244078 237396 244258 237484
rect 244366 237396 244546 237484
rect 244654 237396 244834 237484
rect 244942 237396 245122 237484
rect 245230 237396 245410 237484
rect 245664 237396 245844 237484
rect 245952 237396 246132 237484
rect 246240 237396 246420 237484
rect 246528 237396 246708 237484
rect 246816 237396 246996 237484
rect 247104 237396 247284 237484
rect 247392 237396 247572 237484
rect 247680 237396 247860 237484
rect 248114 237396 248294 237484
rect 248402 237396 248582 237484
rect 248690 237396 248870 237484
rect 248978 237396 249158 237484
rect 249266 237396 249446 237484
rect 249554 237396 249734 237484
rect 249842 237396 250022 237484
rect 250130 237396 250310 237484
rect 250564 237396 250744 237484
rect 360436 237396 360560 237484
rect 360814 237396 360994 237484
rect 361102 237396 361282 237484
rect 361390 237396 361570 237484
rect 361678 237396 361858 237484
rect 361966 237396 362146 237484
rect 362254 237396 362434 237484
rect 362542 237396 362722 237484
rect 362830 237396 363010 237484
rect 363264 237396 363444 237484
rect 363552 237396 363732 237484
rect 363840 237396 364020 237484
rect 364128 237396 364308 237484
rect 364416 237396 364596 237484
rect 364704 237396 364884 237484
rect 364992 237396 365172 237484
rect 365280 237396 365460 237484
rect 365714 237396 365894 237484
rect 366002 237396 366182 237484
rect 366290 237396 366470 237484
rect 366578 237396 366758 237484
rect 366866 237396 367046 237484
rect 367154 237396 367334 237484
rect 367442 237396 367622 237484
rect 367730 237396 367910 237484
rect 243214 237180 243394 237268
rect 243502 237180 243682 237268
rect 243790 237180 243970 237268
rect 244078 237180 244258 237268
rect 244366 237180 244546 237268
rect 244654 237180 244834 237268
rect 244942 237180 245122 237268
rect 245230 237180 245410 237268
rect 245664 237180 245844 237268
rect 245952 237180 246132 237268
rect 246240 237180 246420 237268
rect 246528 237180 246708 237268
rect 246816 237180 246996 237268
rect 247104 237180 247284 237268
rect 247392 237180 247572 237268
rect 247680 237180 247860 237268
rect 248114 237180 248294 237268
rect 248402 237180 248582 237268
rect 248690 237180 248870 237268
rect 248978 237180 249158 237268
rect 249266 237180 249446 237268
rect 249554 237180 249734 237268
rect 249842 237180 250022 237268
rect 250130 237180 250310 237268
rect 250564 237180 250744 237268
rect 360436 237180 360560 237268
rect 360814 237180 360994 237268
rect 361102 237180 361282 237268
rect 361390 237180 361570 237268
rect 361678 237180 361858 237268
rect 361966 237180 362146 237268
rect 362254 237180 362434 237268
rect 362542 237180 362722 237268
rect 362830 237180 363010 237268
rect 363264 237180 363444 237268
rect 363552 237180 363732 237268
rect 363840 237180 364020 237268
rect 364128 237180 364308 237268
rect 364416 237180 364596 237268
rect 364704 237180 364884 237268
rect 364992 237180 365172 237268
rect 365280 237180 365460 237268
rect 365714 237180 365894 237268
rect 366002 237180 366182 237268
rect 366290 237180 366470 237268
rect 366578 237180 366758 237268
rect 366866 237180 367046 237268
rect 367154 237180 367334 237268
rect 367442 237180 367622 237268
rect 367730 237180 367910 237268
rect 243214 236704 243394 236792
rect 243502 236704 243682 236792
rect 243790 236704 243970 236792
rect 244078 236704 244258 236792
rect 244366 236704 244546 236792
rect 244654 236704 244834 236792
rect 244942 236704 245122 236792
rect 245230 236704 245410 236792
rect 245664 236704 245844 236792
rect 245952 236704 246132 236792
rect 246240 236704 246420 236792
rect 246528 236704 246708 236792
rect 246816 236704 246996 236792
rect 247104 236704 247284 236792
rect 247392 236704 247572 236792
rect 247680 236704 247860 236792
rect 248114 236704 248294 236792
rect 248402 236704 248582 236792
rect 248690 236704 248870 236792
rect 248978 236704 249158 236792
rect 249266 236704 249446 236792
rect 249554 236704 249734 236792
rect 249842 236704 250022 236792
rect 250130 236704 250310 236792
rect 250564 236704 250744 236792
rect 360436 236704 360560 236792
rect 360814 236704 360994 236792
rect 361102 236704 361282 236792
rect 361390 236704 361570 236792
rect 361678 236704 361858 236792
rect 361966 236704 362146 236792
rect 362254 236704 362434 236792
rect 362542 236704 362722 236792
rect 362830 236704 363010 236792
rect 363264 236704 363444 236792
rect 363552 236704 363732 236792
rect 363840 236704 364020 236792
rect 364128 236704 364308 236792
rect 364416 236704 364596 236792
rect 364704 236704 364884 236792
rect 364992 236704 365172 236792
rect 365280 236704 365460 236792
rect 365714 236704 365894 236792
rect 366002 236704 366182 236792
rect 366290 236704 366470 236792
rect 366578 236704 366758 236792
rect 366866 236704 367046 236792
rect 367154 236704 367334 236792
rect 367442 236704 367622 236792
rect 367730 236704 367910 236792
rect 243214 236230 243394 236318
rect 243502 236230 243682 236318
rect 243790 236230 243970 236318
rect 244078 236230 244258 236318
rect 244366 236230 244546 236318
rect 244654 236230 244834 236318
rect 244942 236230 245122 236318
rect 245230 236230 245410 236318
rect 245664 236230 245844 236318
rect 245952 236230 246132 236318
rect 246240 236230 246420 236318
rect 246528 236230 246708 236318
rect 246816 236230 246996 236318
rect 247104 236230 247284 236318
rect 247392 236230 247572 236318
rect 247680 236230 247860 236318
rect 248114 236230 248294 236318
rect 248402 236230 248582 236318
rect 248690 236230 248870 236318
rect 248978 236230 249158 236318
rect 249266 236230 249446 236318
rect 249554 236230 249734 236318
rect 249842 236230 250022 236318
rect 250130 236230 250310 236318
rect 250564 236230 250744 236318
rect 360436 236230 360560 236318
rect 360814 236230 360994 236318
rect 361102 236230 361282 236318
rect 361390 236230 361570 236318
rect 361678 236230 361858 236318
rect 361966 236230 362146 236318
rect 362254 236230 362434 236318
rect 362542 236230 362722 236318
rect 362830 236230 363010 236318
rect 363264 236230 363444 236318
rect 363552 236230 363732 236318
rect 363840 236230 364020 236318
rect 364128 236230 364308 236318
rect 364416 236230 364596 236318
rect 364704 236230 364884 236318
rect 364992 236230 365172 236318
rect 365280 236230 365460 236318
rect 365714 236230 365894 236318
rect 366002 236230 366182 236318
rect 366290 236230 366470 236318
rect 366578 236230 366758 236318
rect 366866 236230 367046 236318
rect 367154 236230 367334 236318
rect 367442 236230 367622 236318
rect 367730 236230 367910 236318
rect 243214 235754 243394 235842
rect 243502 235754 243682 235842
rect 243790 235754 243970 235842
rect 244078 235754 244258 235842
rect 244366 235754 244546 235842
rect 244654 235754 244834 235842
rect 244942 235754 245122 235842
rect 245230 235754 245410 235842
rect 245664 235754 245844 235842
rect 245952 235754 246132 235842
rect 246240 235754 246420 235842
rect 246528 235754 246708 235842
rect 246816 235754 246996 235842
rect 247104 235754 247284 235842
rect 247392 235754 247572 235842
rect 247680 235754 247860 235842
rect 248114 235754 248294 235842
rect 248402 235754 248582 235842
rect 248690 235754 248870 235842
rect 248978 235754 249158 235842
rect 249266 235754 249446 235842
rect 249554 235754 249734 235842
rect 249842 235754 250022 235842
rect 250130 235754 250310 235842
rect 250564 235754 250744 235842
rect 360436 235754 360560 235842
rect 360814 235754 360994 235842
rect 361102 235754 361282 235842
rect 361390 235754 361570 235842
rect 361678 235754 361858 235842
rect 361966 235754 362146 235842
rect 362254 235754 362434 235842
rect 362542 235754 362722 235842
rect 362830 235754 363010 235842
rect 363264 235754 363444 235842
rect 363552 235754 363732 235842
rect 363840 235754 364020 235842
rect 364128 235754 364308 235842
rect 364416 235754 364596 235842
rect 364704 235754 364884 235842
rect 364992 235754 365172 235842
rect 365280 235754 365460 235842
rect 365714 235754 365894 235842
rect 366002 235754 366182 235842
rect 366290 235754 366470 235842
rect 366578 235754 366758 235842
rect 366866 235754 367046 235842
rect 367154 235754 367334 235842
rect 367442 235754 367622 235842
rect 367730 235754 367910 235842
rect 243214 235538 243394 235626
rect 243502 235538 243682 235626
rect 243790 235538 243970 235626
rect 244078 235538 244258 235626
rect 244366 235538 244546 235626
rect 244654 235538 244834 235626
rect 244942 235538 245122 235626
rect 245230 235538 245410 235626
rect 245664 235538 245844 235626
rect 245952 235538 246132 235626
rect 246240 235538 246420 235626
rect 246528 235538 246708 235626
rect 246816 235538 246996 235626
rect 247104 235538 247284 235626
rect 247392 235538 247572 235626
rect 247680 235538 247860 235626
rect 248114 235538 248294 235626
rect 248402 235538 248582 235626
rect 248690 235538 248870 235626
rect 248978 235538 249158 235626
rect 249266 235538 249446 235626
rect 249554 235538 249734 235626
rect 249842 235538 250022 235626
rect 250130 235538 250310 235626
rect 250564 235538 250744 235626
rect 360436 235538 360560 235626
rect 360814 235538 360994 235626
rect 361102 235538 361282 235626
rect 361390 235538 361570 235626
rect 361678 235538 361858 235626
rect 361966 235538 362146 235626
rect 362254 235538 362434 235626
rect 362542 235538 362722 235626
rect 362830 235538 363010 235626
rect 363264 235538 363444 235626
rect 363552 235538 363732 235626
rect 363840 235538 364020 235626
rect 364128 235538 364308 235626
rect 364416 235538 364596 235626
rect 364704 235538 364884 235626
rect 364992 235538 365172 235626
rect 365280 235538 365460 235626
rect 365714 235538 365894 235626
rect 366002 235538 366182 235626
rect 366290 235538 366470 235626
rect 366578 235538 366758 235626
rect 366866 235538 367046 235626
rect 367154 235538 367334 235626
rect 367442 235538 367622 235626
rect 367730 235538 367910 235626
rect 243214 235062 243394 235150
rect 243502 235062 243682 235150
rect 243790 235062 243970 235150
rect 244078 235062 244258 235150
rect 244366 235062 244546 235150
rect 244654 235062 244834 235150
rect 244942 235062 245122 235150
rect 245230 235062 245410 235150
rect 245664 235062 245844 235150
rect 245952 235062 246132 235150
rect 246240 235062 246420 235150
rect 246528 235062 246708 235150
rect 246816 235062 246996 235150
rect 247104 235062 247284 235150
rect 247392 235062 247572 235150
rect 247680 235062 247860 235150
rect 248114 235062 248294 235150
rect 248402 235062 248582 235150
rect 248690 235062 248870 235150
rect 248978 235062 249158 235150
rect 249266 235062 249446 235150
rect 249554 235062 249734 235150
rect 249842 235062 250022 235150
rect 250130 235062 250310 235150
rect 250564 235062 250744 235150
rect 360436 235062 360560 235150
rect 360814 235062 360994 235150
rect 361102 235062 361282 235150
rect 361390 235062 361570 235150
rect 361678 235062 361858 235150
rect 361966 235062 362146 235150
rect 362254 235062 362434 235150
rect 362542 235062 362722 235150
rect 362830 235062 363010 235150
rect 363264 235062 363444 235150
rect 363552 235062 363732 235150
rect 363840 235062 364020 235150
rect 364128 235062 364308 235150
rect 364416 235062 364596 235150
rect 364704 235062 364884 235150
rect 364992 235062 365172 235150
rect 365280 235062 365460 235150
rect 365714 235062 365894 235150
rect 366002 235062 366182 235150
rect 366290 235062 366470 235150
rect 366578 235062 366758 235150
rect 366866 235062 367046 235150
rect 367154 235062 367334 235150
rect 367442 235062 367622 235150
rect 367730 235062 367910 235150
rect 243214 234846 243394 234934
rect 243502 234846 243682 234934
rect 243790 234846 243970 234934
rect 244078 234846 244258 234934
rect 244366 234846 244546 234934
rect 244654 234846 244834 234934
rect 244942 234846 245122 234934
rect 245230 234846 245410 234934
rect 245664 234846 245844 234934
rect 245952 234846 246132 234934
rect 246240 234846 246420 234934
rect 246528 234846 246708 234934
rect 246816 234846 246996 234934
rect 247104 234846 247284 234934
rect 247392 234846 247572 234934
rect 247680 234846 247860 234934
rect 248114 234846 248294 234934
rect 248402 234846 248582 234934
rect 248690 234846 248870 234934
rect 248978 234846 249158 234934
rect 249266 234846 249446 234934
rect 249554 234846 249734 234934
rect 249842 234846 250022 234934
rect 250130 234846 250310 234934
rect 250564 234846 250744 234934
rect 360436 234846 360560 234934
rect 360814 234846 360994 234934
rect 361102 234846 361282 234934
rect 361390 234846 361570 234934
rect 361678 234846 361858 234934
rect 361966 234846 362146 234934
rect 362254 234846 362434 234934
rect 362542 234846 362722 234934
rect 362830 234846 363010 234934
rect 363264 234846 363444 234934
rect 363552 234846 363732 234934
rect 363840 234846 364020 234934
rect 364128 234846 364308 234934
rect 364416 234846 364596 234934
rect 364704 234846 364884 234934
rect 364992 234846 365172 234934
rect 365280 234846 365460 234934
rect 365714 234846 365894 234934
rect 366002 234846 366182 234934
rect 366290 234846 366470 234934
rect 366578 234846 366758 234934
rect 366866 234846 367046 234934
rect 367154 234846 367334 234934
rect 367442 234846 367622 234934
rect 367730 234846 367910 234934
rect 243214 234370 243394 234458
rect 243502 234370 243682 234458
rect 243790 234370 243970 234458
rect 244078 234370 244258 234458
rect 244366 234370 244546 234458
rect 244654 234370 244834 234458
rect 244942 234370 245122 234458
rect 245230 234370 245410 234458
rect 245664 234370 245844 234458
rect 245952 234370 246132 234458
rect 246240 234370 246420 234458
rect 246528 234370 246708 234458
rect 246816 234370 246996 234458
rect 247104 234370 247284 234458
rect 247392 234370 247572 234458
rect 247680 234370 247860 234458
rect 248114 234370 248294 234458
rect 248402 234370 248582 234458
rect 248690 234370 248870 234458
rect 248978 234370 249158 234458
rect 249266 234370 249446 234458
rect 249554 234370 249734 234458
rect 249842 234370 250022 234458
rect 250130 234370 250310 234458
rect 250564 234370 250744 234458
rect 360436 234370 360560 234458
rect 360814 234370 360994 234458
rect 361102 234370 361282 234458
rect 361390 234370 361570 234458
rect 361678 234370 361858 234458
rect 361966 234370 362146 234458
rect 362254 234370 362434 234458
rect 362542 234370 362722 234458
rect 362830 234370 363010 234458
rect 363264 234370 363444 234458
rect 363552 234370 363732 234458
rect 363840 234370 364020 234458
rect 364128 234370 364308 234458
rect 364416 234370 364596 234458
rect 364704 234370 364884 234458
rect 364992 234370 365172 234458
rect 365280 234370 365460 234458
rect 365714 234370 365894 234458
rect 366002 234370 366182 234458
rect 366290 234370 366470 234458
rect 366578 234370 366758 234458
rect 366866 234370 367046 234458
rect 367154 234370 367334 234458
rect 367442 234370 367622 234458
rect 367730 234370 367910 234458
rect 243214 234154 243394 234242
rect 243502 234154 243682 234242
rect 243790 234154 243970 234242
rect 244078 234154 244258 234242
rect 244366 234154 244546 234242
rect 244654 234154 244834 234242
rect 244942 234154 245122 234242
rect 245230 234154 245410 234242
rect 245664 234154 245844 234242
rect 245952 234154 246132 234242
rect 246240 234154 246420 234242
rect 246528 234154 246708 234242
rect 246816 234154 246996 234242
rect 247104 234154 247284 234242
rect 247392 234154 247572 234242
rect 247680 234154 247860 234242
rect 248114 234154 248294 234242
rect 248402 234154 248582 234242
rect 248690 234154 248870 234242
rect 248978 234154 249158 234242
rect 249266 234154 249446 234242
rect 249554 234154 249734 234242
rect 249842 234154 250022 234242
rect 250130 234154 250310 234242
rect 250564 234154 250744 234242
rect 360436 234154 360560 234242
rect 360814 234154 360994 234242
rect 361102 234154 361282 234242
rect 361390 234154 361570 234242
rect 361678 234154 361858 234242
rect 361966 234154 362146 234242
rect 362254 234154 362434 234242
rect 362542 234154 362722 234242
rect 362830 234154 363010 234242
rect 363264 234154 363444 234242
rect 363552 234154 363732 234242
rect 363840 234154 364020 234242
rect 364128 234154 364308 234242
rect 364416 234154 364596 234242
rect 364704 234154 364884 234242
rect 364992 234154 365172 234242
rect 365280 234154 365460 234242
rect 365714 234154 365894 234242
rect 366002 234154 366182 234242
rect 366290 234154 366470 234242
rect 366578 234154 366758 234242
rect 366866 234154 367046 234242
rect 367154 234154 367334 234242
rect 367442 234154 367622 234242
rect 367730 234154 367910 234242
rect 243214 233678 243394 233766
rect 243502 233678 243682 233766
rect 243790 233678 243970 233766
rect 244078 233678 244258 233766
rect 244366 233678 244546 233766
rect 244654 233678 244834 233766
rect 244942 233678 245122 233766
rect 245230 233678 245410 233766
rect 245664 233678 245844 233766
rect 245952 233678 246132 233766
rect 246240 233678 246420 233766
rect 246528 233678 246708 233766
rect 246816 233678 246996 233766
rect 247104 233678 247284 233766
rect 247392 233678 247572 233766
rect 247680 233678 247860 233766
rect 248114 233678 248294 233766
rect 248402 233678 248582 233766
rect 248690 233678 248870 233766
rect 248978 233678 249158 233766
rect 249266 233678 249446 233766
rect 249554 233678 249734 233766
rect 249842 233678 250022 233766
rect 250130 233678 250310 233766
rect 250564 233678 250744 233766
rect 360436 233678 360560 233766
rect 360814 233678 360994 233766
rect 361102 233678 361282 233766
rect 361390 233678 361570 233766
rect 361678 233678 361858 233766
rect 361966 233678 362146 233766
rect 362254 233678 362434 233766
rect 362542 233678 362722 233766
rect 362830 233678 363010 233766
rect 363264 233678 363444 233766
rect 363552 233678 363732 233766
rect 363840 233678 364020 233766
rect 364128 233678 364308 233766
rect 364416 233678 364596 233766
rect 364704 233678 364884 233766
rect 364992 233678 365172 233766
rect 365280 233678 365460 233766
rect 365714 233678 365894 233766
rect 366002 233678 366182 233766
rect 366290 233678 366470 233766
rect 366578 233678 366758 233766
rect 366866 233678 367046 233766
rect 367154 233678 367334 233766
rect 367442 233678 367622 233766
rect 367730 233678 367910 233766
rect 243214 233204 243394 233292
rect 243502 233204 243682 233292
rect 243790 233204 243970 233292
rect 244078 233204 244258 233292
rect 244366 233204 244546 233292
rect 244654 233204 244834 233292
rect 244942 233204 245122 233292
rect 245230 233204 245410 233292
rect 245664 233204 245844 233292
rect 245952 233204 246132 233292
rect 246240 233204 246420 233292
rect 246528 233204 246708 233292
rect 246816 233204 246996 233292
rect 247104 233204 247284 233292
rect 247392 233204 247572 233292
rect 247680 233204 247860 233292
rect 248114 233204 248294 233292
rect 248402 233204 248582 233292
rect 248690 233204 248870 233292
rect 248978 233204 249158 233292
rect 249266 233204 249446 233292
rect 249554 233204 249734 233292
rect 249842 233204 250022 233292
rect 250130 233204 250310 233292
rect 250564 233204 250744 233292
rect 360436 233204 360560 233292
rect 360814 233204 360994 233292
rect 361102 233204 361282 233292
rect 361390 233204 361570 233292
rect 361678 233204 361858 233292
rect 361966 233204 362146 233292
rect 362254 233204 362434 233292
rect 362542 233204 362722 233292
rect 362830 233204 363010 233292
rect 363264 233204 363444 233292
rect 363552 233204 363732 233292
rect 363840 233204 364020 233292
rect 364128 233204 364308 233292
rect 364416 233204 364596 233292
rect 364704 233204 364884 233292
rect 364992 233204 365172 233292
rect 365280 233204 365460 233292
rect 365714 233204 365894 233292
rect 366002 233204 366182 233292
rect 366290 233204 366470 233292
rect 366578 233204 366758 233292
rect 366866 233204 367046 233292
rect 367154 233204 367334 233292
rect 367442 233204 367622 233292
rect 367730 233204 367910 233292
rect 243214 232728 243394 232816
rect 243502 232728 243682 232816
rect 243790 232728 243970 232816
rect 244078 232728 244258 232816
rect 244366 232728 244546 232816
rect 244654 232728 244834 232816
rect 244942 232728 245122 232816
rect 245230 232728 245410 232816
rect 245664 232728 245844 232816
rect 245952 232728 246132 232816
rect 246240 232728 246420 232816
rect 246528 232728 246708 232816
rect 246816 232728 246996 232816
rect 247104 232728 247284 232816
rect 247392 232728 247572 232816
rect 247680 232728 247860 232816
rect 248114 232728 248294 232816
rect 248402 232728 248582 232816
rect 248690 232728 248870 232816
rect 248978 232728 249158 232816
rect 249266 232728 249446 232816
rect 249554 232728 249734 232816
rect 249842 232728 250022 232816
rect 250130 232728 250310 232816
rect 250564 232728 250744 232816
rect 360436 232728 360560 232816
rect 360814 232728 360994 232816
rect 361102 232728 361282 232816
rect 361390 232728 361570 232816
rect 361678 232728 361858 232816
rect 361966 232728 362146 232816
rect 362254 232728 362434 232816
rect 362542 232728 362722 232816
rect 362830 232728 363010 232816
rect 363264 232728 363444 232816
rect 363552 232728 363732 232816
rect 363840 232728 364020 232816
rect 364128 232728 364308 232816
rect 364416 232728 364596 232816
rect 364704 232728 364884 232816
rect 364992 232728 365172 232816
rect 365280 232728 365460 232816
rect 365714 232728 365894 232816
rect 366002 232728 366182 232816
rect 366290 232728 366470 232816
rect 366578 232728 366758 232816
rect 366866 232728 367046 232816
rect 367154 232728 367334 232816
rect 367442 232728 367622 232816
rect 367730 232728 367910 232816
rect 243214 232512 243394 232600
rect 243502 232512 243682 232600
rect 243790 232512 243970 232600
rect 244078 232512 244258 232600
rect 244366 232512 244546 232600
rect 244654 232512 244834 232600
rect 244942 232512 245122 232600
rect 245230 232512 245410 232600
rect 245664 232512 245844 232600
rect 245952 232512 246132 232600
rect 246240 232512 246420 232600
rect 246528 232512 246708 232600
rect 246816 232512 246996 232600
rect 247104 232512 247284 232600
rect 247392 232512 247572 232600
rect 247680 232512 247860 232600
rect 248114 232512 248294 232600
rect 248402 232512 248582 232600
rect 248690 232512 248870 232600
rect 248978 232512 249158 232600
rect 249266 232512 249446 232600
rect 249554 232512 249734 232600
rect 249842 232512 250022 232600
rect 250130 232512 250310 232600
rect 250564 232512 250744 232600
rect 360436 232512 360560 232600
rect 360814 232512 360994 232600
rect 361102 232512 361282 232600
rect 361390 232512 361570 232600
rect 361678 232512 361858 232600
rect 361966 232512 362146 232600
rect 362254 232512 362434 232600
rect 362542 232512 362722 232600
rect 362830 232512 363010 232600
rect 363264 232512 363444 232600
rect 363552 232512 363732 232600
rect 363840 232512 364020 232600
rect 364128 232512 364308 232600
rect 364416 232512 364596 232600
rect 364704 232512 364884 232600
rect 364992 232512 365172 232600
rect 365280 232512 365460 232600
rect 365714 232512 365894 232600
rect 366002 232512 366182 232600
rect 366290 232512 366470 232600
rect 366578 232512 366758 232600
rect 366866 232512 367046 232600
rect 367154 232512 367334 232600
rect 367442 232512 367622 232600
rect 367730 232512 367910 232600
rect 243214 232036 243394 232124
rect 243502 232036 243682 232124
rect 243790 232036 243970 232124
rect 244078 232036 244258 232124
rect 244366 232036 244546 232124
rect 244654 232036 244834 232124
rect 244942 232036 245122 232124
rect 245230 232036 245410 232124
rect 245664 232036 245844 232124
rect 245952 232036 246132 232124
rect 246240 232036 246420 232124
rect 246528 232036 246708 232124
rect 246816 232036 246996 232124
rect 247104 232036 247284 232124
rect 247392 232036 247572 232124
rect 247680 232036 247860 232124
rect 248114 232036 248294 232124
rect 248402 232036 248582 232124
rect 248690 232036 248870 232124
rect 248978 232036 249158 232124
rect 249266 232036 249446 232124
rect 249554 232036 249734 232124
rect 249842 232036 250022 232124
rect 250130 232036 250310 232124
rect 250564 232036 250744 232124
rect 360436 232036 360560 232124
rect 360814 232036 360994 232124
rect 361102 232036 361282 232124
rect 361390 232036 361570 232124
rect 361678 232036 361858 232124
rect 361966 232036 362146 232124
rect 362254 232036 362434 232124
rect 362542 232036 362722 232124
rect 362830 232036 363010 232124
rect 363264 232036 363444 232124
rect 363552 232036 363732 232124
rect 363840 232036 364020 232124
rect 364128 232036 364308 232124
rect 364416 232036 364596 232124
rect 364704 232036 364884 232124
rect 364992 232036 365172 232124
rect 365280 232036 365460 232124
rect 365714 232036 365894 232124
rect 366002 232036 366182 232124
rect 366290 232036 366470 232124
rect 366578 232036 366758 232124
rect 366866 232036 367046 232124
rect 367154 232036 367334 232124
rect 367442 232036 367622 232124
rect 367730 232036 367910 232124
rect 243214 231820 243394 231908
rect 243502 231820 243682 231908
rect 243790 231820 243970 231908
rect 244078 231820 244258 231908
rect 244366 231820 244546 231908
rect 244654 231820 244834 231908
rect 244942 231820 245122 231908
rect 245230 231820 245410 231908
rect 245664 231820 245844 231908
rect 245952 231820 246132 231908
rect 246240 231820 246420 231908
rect 246528 231820 246708 231908
rect 246816 231820 246996 231908
rect 247104 231820 247284 231908
rect 247392 231820 247572 231908
rect 247680 231820 247860 231908
rect 248114 231820 248294 231908
rect 248402 231820 248582 231908
rect 248690 231820 248870 231908
rect 248978 231820 249158 231908
rect 249266 231820 249446 231908
rect 249554 231820 249734 231908
rect 249842 231820 250022 231908
rect 250130 231820 250310 231908
rect 250564 231820 250744 231908
rect 360436 231820 360560 231908
rect 360814 231820 360994 231908
rect 361102 231820 361282 231908
rect 361390 231820 361570 231908
rect 361678 231820 361858 231908
rect 361966 231820 362146 231908
rect 362254 231820 362434 231908
rect 362542 231820 362722 231908
rect 362830 231820 363010 231908
rect 363264 231820 363444 231908
rect 363552 231820 363732 231908
rect 363840 231820 364020 231908
rect 364128 231820 364308 231908
rect 364416 231820 364596 231908
rect 364704 231820 364884 231908
rect 364992 231820 365172 231908
rect 365280 231820 365460 231908
rect 365714 231820 365894 231908
rect 366002 231820 366182 231908
rect 366290 231820 366470 231908
rect 366578 231820 366758 231908
rect 366866 231820 367046 231908
rect 367154 231820 367334 231908
rect 367442 231820 367622 231908
rect 367730 231820 367910 231908
rect 243214 231344 243394 231432
rect 243502 231344 243682 231432
rect 243790 231344 243970 231432
rect 244078 231344 244258 231432
rect 244366 231344 244546 231432
rect 244654 231344 244834 231432
rect 244942 231344 245122 231432
rect 245230 231344 245410 231432
rect 245664 231344 245844 231432
rect 245952 231344 246132 231432
rect 246240 231344 246420 231432
rect 246528 231344 246708 231432
rect 246816 231344 246996 231432
rect 247104 231344 247284 231432
rect 247392 231344 247572 231432
rect 247680 231344 247860 231432
rect 248114 231344 248294 231432
rect 248402 231344 248582 231432
rect 248690 231344 248870 231432
rect 248978 231344 249158 231432
rect 249266 231344 249446 231432
rect 249554 231344 249734 231432
rect 249842 231344 250022 231432
rect 250130 231344 250310 231432
rect 250564 231344 250744 231432
rect 360436 231344 360560 231432
rect 360814 231344 360994 231432
rect 361102 231344 361282 231432
rect 361390 231344 361570 231432
rect 361678 231344 361858 231432
rect 361966 231344 362146 231432
rect 362254 231344 362434 231432
rect 362542 231344 362722 231432
rect 362830 231344 363010 231432
rect 363264 231344 363444 231432
rect 363552 231344 363732 231432
rect 363840 231344 364020 231432
rect 364128 231344 364308 231432
rect 364416 231344 364596 231432
rect 364704 231344 364884 231432
rect 364992 231344 365172 231432
rect 365280 231344 365460 231432
rect 365714 231344 365894 231432
rect 366002 231344 366182 231432
rect 366290 231344 366470 231432
rect 366578 231344 366758 231432
rect 366866 231344 367046 231432
rect 367154 231344 367334 231432
rect 367442 231344 367622 231432
rect 367730 231344 367910 231432
rect 243214 231128 243394 231216
rect 243502 231128 243682 231216
rect 243790 231128 243970 231216
rect 244078 231128 244258 231216
rect 244366 231128 244546 231216
rect 244654 231128 244834 231216
rect 244942 231128 245122 231216
rect 245230 231128 245410 231216
rect 245664 231128 245844 231216
rect 245952 231128 246132 231216
rect 246240 231128 246420 231216
rect 246528 231128 246708 231216
rect 246816 231128 246996 231216
rect 247104 231128 247284 231216
rect 247392 231128 247572 231216
rect 247680 231128 247860 231216
rect 248114 231128 248294 231216
rect 248402 231128 248582 231216
rect 248690 231128 248870 231216
rect 248978 231128 249158 231216
rect 249266 231128 249446 231216
rect 249554 231128 249734 231216
rect 249842 231128 250022 231216
rect 250130 231128 250310 231216
rect 250564 231128 250744 231216
rect 360436 231128 360560 231216
rect 360814 231128 360994 231216
rect 361102 231128 361282 231216
rect 361390 231128 361570 231216
rect 361678 231128 361858 231216
rect 361966 231128 362146 231216
rect 362254 231128 362434 231216
rect 362542 231128 362722 231216
rect 362830 231128 363010 231216
rect 363264 231128 363444 231216
rect 363552 231128 363732 231216
rect 363840 231128 364020 231216
rect 364128 231128 364308 231216
rect 364416 231128 364596 231216
rect 364704 231128 364884 231216
rect 364992 231128 365172 231216
rect 365280 231128 365460 231216
rect 365714 231128 365894 231216
rect 366002 231128 366182 231216
rect 366290 231128 366470 231216
rect 366578 231128 366758 231216
rect 366866 231128 367046 231216
rect 367154 231128 367334 231216
rect 367442 231128 367622 231216
rect 367730 231128 367910 231216
rect 243214 230652 243394 230740
rect 243502 230652 243682 230740
rect 243790 230652 243970 230740
rect 244078 230652 244258 230740
rect 244366 230652 244546 230740
rect 244654 230652 244834 230740
rect 244942 230652 245122 230740
rect 245230 230652 245410 230740
rect 245664 230652 245844 230740
rect 245952 230652 246132 230740
rect 246240 230652 246420 230740
rect 246528 230652 246708 230740
rect 246816 230652 246996 230740
rect 247104 230652 247284 230740
rect 247392 230652 247572 230740
rect 247680 230652 247860 230740
rect 248114 230652 248294 230740
rect 248402 230652 248582 230740
rect 248690 230652 248870 230740
rect 248978 230652 249158 230740
rect 249266 230652 249446 230740
rect 249554 230652 249734 230740
rect 249842 230652 250022 230740
rect 250130 230652 250310 230740
rect 250564 230652 250744 230740
rect 360436 230652 360560 230740
rect 360814 230652 360994 230740
rect 361102 230652 361282 230740
rect 361390 230652 361570 230740
rect 361678 230652 361858 230740
rect 361966 230652 362146 230740
rect 362254 230652 362434 230740
rect 362542 230652 362722 230740
rect 362830 230652 363010 230740
rect 363264 230652 363444 230740
rect 363552 230652 363732 230740
rect 363840 230652 364020 230740
rect 364128 230652 364308 230740
rect 364416 230652 364596 230740
rect 364704 230652 364884 230740
rect 364992 230652 365172 230740
rect 365280 230652 365460 230740
rect 365714 230652 365894 230740
rect 366002 230652 366182 230740
rect 366290 230652 366470 230740
rect 366578 230652 366758 230740
rect 366866 230652 367046 230740
rect 367154 230652 367334 230740
rect 367442 230652 367622 230740
rect 367730 230652 367910 230740
rect 243214 230178 243394 230266
rect 243502 230178 243682 230266
rect 243790 230178 243970 230266
rect 244078 230178 244258 230266
rect 244366 230178 244546 230266
rect 244654 230178 244834 230266
rect 244942 230178 245122 230266
rect 245230 230178 245410 230266
rect 245664 230178 245844 230266
rect 245952 230178 246132 230266
rect 246240 230178 246420 230266
rect 246528 230178 246708 230266
rect 246816 230178 246996 230266
rect 247104 230178 247284 230266
rect 247392 230178 247572 230266
rect 247680 230178 247860 230266
rect 248114 230178 248294 230266
rect 248402 230178 248582 230266
rect 248690 230178 248870 230266
rect 248978 230178 249158 230266
rect 249266 230178 249446 230266
rect 249554 230178 249734 230266
rect 249842 230178 250022 230266
rect 250130 230178 250310 230266
rect 250564 230178 250744 230266
rect 360436 230178 360560 230266
rect 360814 230178 360994 230266
rect 361102 230178 361282 230266
rect 361390 230178 361570 230266
rect 361678 230178 361858 230266
rect 361966 230178 362146 230266
rect 362254 230178 362434 230266
rect 362542 230178 362722 230266
rect 362830 230178 363010 230266
rect 363264 230178 363444 230266
rect 363552 230178 363732 230266
rect 363840 230178 364020 230266
rect 364128 230178 364308 230266
rect 364416 230178 364596 230266
rect 364704 230178 364884 230266
rect 364992 230178 365172 230266
rect 365280 230178 365460 230266
rect 365714 230178 365894 230266
rect 366002 230178 366182 230266
rect 366290 230178 366470 230266
rect 366578 230178 366758 230266
rect 366866 230178 367046 230266
rect 367154 230178 367334 230266
rect 367442 230178 367622 230266
rect 367730 230178 367910 230266
rect 243214 229702 243394 229790
rect 243502 229702 243682 229790
rect 243790 229702 243970 229790
rect 244078 229702 244258 229790
rect 244366 229702 244546 229790
rect 244654 229702 244834 229790
rect 244942 229702 245122 229790
rect 245230 229702 245410 229790
rect 245664 229702 245844 229790
rect 245952 229702 246132 229790
rect 246240 229702 246420 229790
rect 246528 229702 246708 229790
rect 246816 229702 246996 229790
rect 247104 229702 247284 229790
rect 247392 229702 247572 229790
rect 247680 229702 247860 229790
rect 248114 229702 248294 229790
rect 248402 229702 248582 229790
rect 248690 229702 248870 229790
rect 248978 229702 249158 229790
rect 249266 229702 249446 229790
rect 249554 229702 249734 229790
rect 249842 229702 250022 229790
rect 250130 229702 250310 229790
rect 250564 229702 250744 229790
rect 360436 229702 360560 229790
rect 360814 229702 360994 229790
rect 361102 229702 361282 229790
rect 361390 229702 361570 229790
rect 361678 229702 361858 229790
rect 361966 229702 362146 229790
rect 362254 229702 362434 229790
rect 362542 229702 362722 229790
rect 362830 229702 363010 229790
rect 363264 229702 363444 229790
rect 363552 229702 363732 229790
rect 363840 229702 364020 229790
rect 364128 229702 364308 229790
rect 364416 229702 364596 229790
rect 364704 229702 364884 229790
rect 364992 229702 365172 229790
rect 365280 229702 365460 229790
rect 365714 229702 365894 229790
rect 366002 229702 366182 229790
rect 366290 229702 366470 229790
rect 366578 229702 366758 229790
rect 366866 229702 367046 229790
rect 367154 229702 367334 229790
rect 367442 229702 367622 229790
rect 367730 229702 367910 229790
rect 243214 229486 243394 229574
rect 243502 229486 243682 229574
rect 243790 229486 243970 229574
rect 244078 229486 244258 229574
rect 244366 229486 244546 229574
rect 244654 229486 244834 229574
rect 244942 229486 245122 229574
rect 245230 229486 245410 229574
rect 245664 229486 245844 229574
rect 245952 229486 246132 229574
rect 246240 229486 246420 229574
rect 246528 229486 246708 229574
rect 246816 229486 246996 229574
rect 247104 229486 247284 229574
rect 247392 229486 247572 229574
rect 247680 229486 247860 229574
rect 248114 229486 248294 229574
rect 248402 229486 248582 229574
rect 248690 229486 248870 229574
rect 248978 229486 249158 229574
rect 249266 229486 249446 229574
rect 249554 229486 249734 229574
rect 249842 229486 250022 229574
rect 250130 229486 250310 229574
rect 250564 229486 250744 229574
rect 360436 229486 360560 229574
rect 360814 229486 360994 229574
rect 361102 229486 361282 229574
rect 361390 229486 361570 229574
rect 361678 229486 361858 229574
rect 361966 229486 362146 229574
rect 362254 229486 362434 229574
rect 362542 229486 362722 229574
rect 362830 229486 363010 229574
rect 363264 229486 363444 229574
rect 363552 229486 363732 229574
rect 363840 229486 364020 229574
rect 364128 229486 364308 229574
rect 364416 229486 364596 229574
rect 364704 229486 364884 229574
rect 364992 229486 365172 229574
rect 365280 229486 365460 229574
rect 365714 229486 365894 229574
rect 366002 229486 366182 229574
rect 366290 229486 366470 229574
rect 366578 229486 366758 229574
rect 366866 229486 367046 229574
rect 367154 229486 367334 229574
rect 367442 229486 367622 229574
rect 367730 229486 367910 229574
rect 243214 229010 243394 229098
rect 243502 229010 243682 229098
rect 243790 229010 243970 229098
rect 244078 229010 244258 229098
rect 244366 229010 244546 229098
rect 244654 229010 244834 229098
rect 244942 229010 245122 229098
rect 245230 229010 245410 229098
rect 245664 229010 245844 229098
rect 245952 229010 246132 229098
rect 246240 229010 246420 229098
rect 246528 229010 246708 229098
rect 246816 229010 246996 229098
rect 247104 229010 247284 229098
rect 247392 229010 247572 229098
rect 247680 229010 247860 229098
rect 248114 229010 248294 229098
rect 248402 229010 248582 229098
rect 248690 229010 248870 229098
rect 248978 229010 249158 229098
rect 249266 229010 249446 229098
rect 249554 229010 249734 229098
rect 249842 229010 250022 229098
rect 250130 229010 250310 229098
rect 250564 229010 250744 229098
rect 360436 229010 360560 229098
rect 360814 229010 360994 229098
rect 361102 229010 361282 229098
rect 361390 229010 361570 229098
rect 361678 229010 361858 229098
rect 361966 229010 362146 229098
rect 362254 229010 362434 229098
rect 362542 229010 362722 229098
rect 362830 229010 363010 229098
rect 363264 229010 363444 229098
rect 363552 229010 363732 229098
rect 363840 229010 364020 229098
rect 364128 229010 364308 229098
rect 364416 229010 364596 229098
rect 364704 229010 364884 229098
rect 364992 229010 365172 229098
rect 365280 229010 365460 229098
rect 365714 229010 365894 229098
rect 366002 229010 366182 229098
rect 366290 229010 366470 229098
rect 366578 229010 366758 229098
rect 366866 229010 367046 229098
rect 367154 229010 367334 229098
rect 367442 229010 367622 229098
rect 367730 229010 367910 229098
rect 243214 228794 243394 228882
rect 243502 228794 243682 228882
rect 243790 228794 243970 228882
rect 244078 228794 244258 228882
rect 244366 228794 244546 228882
rect 244654 228794 244834 228882
rect 244942 228794 245122 228882
rect 245230 228794 245410 228882
rect 245664 228794 245844 228882
rect 245952 228794 246132 228882
rect 246240 228794 246420 228882
rect 246528 228794 246708 228882
rect 246816 228794 246996 228882
rect 247104 228794 247284 228882
rect 247392 228794 247572 228882
rect 247680 228794 247860 228882
rect 248114 228794 248294 228882
rect 248402 228794 248582 228882
rect 248690 228794 248870 228882
rect 248978 228794 249158 228882
rect 249266 228794 249446 228882
rect 249554 228794 249734 228882
rect 249842 228794 250022 228882
rect 250130 228794 250310 228882
rect 250564 228794 250744 228882
rect 360436 228794 360560 228882
rect 360814 228794 360994 228882
rect 361102 228794 361282 228882
rect 361390 228794 361570 228882
rect 361678 228794 361858 228882
rect 361966 228794 362146 228882
rect 362254 228794 362434 228882
rect 362542 228794 362722 228882
rect 362830 228794 363010 228882
rect 363264 228794 363444 228882
rect 363552 228794 363732 228882
rect 363840 228794 364020 228882
rect 364128 228794 364308 228882
rect 364416 228794 364596 228882
rect 364704 228794 364884 228882
rect 364992 228794 365172 228882
rect 365280 228794 365460 228882
rect 365714 228794 365894 228882
rect 366002 228794 366182 228882
rect 366290 228794 366470 228882
rect 366578 228794 366758 228882
rect 366866 228794 367046 228882
rect 367154 228794 367334 228882
rect 367442 228794 367622 228882
rect 367730 228794 367910 228882
rect 243214 228318 243394 228406
rect 243502 228318 243682 228406
rect 243790 228318 243970 228406
rect 244078 228318 244258 228406
rect 244366 228318 244546 228406
rect 244654 228318 244834 228406
rect 244942 228318 245122 228406
rect 245230 228318 245410 228406
rect 245664 228318 245844 228406
rect 245952 228318 246132 228406
rect 246240 228318 246420 228406
rect 246528 228318 246708 228406
rect 246816 228318 246996 228406
rect 247104 228318 247284 228406
rect 247392 228318 247572 228406
rect 247680 228318 247860 228406
rect 248114 228318 248294 228406
rect 248402 228318 248582 228406
rect 248690 228318 248870 228406
rect 248978 228318 249158 228406
rect 249266 228318 249446 228406
rect 249554 228318 249734 228406
rect 249842 228318 250022 228406
rect 250130 228318 250310 228406
rect 250564 228318 250744 228406
rect 360436 228318 360560 228406
rect 360814 228318 360994 228406
rect 361102 228318 361282 228406
rect 361390 228318 361570 228406
rect 361678 228318 361858 228406
rect 361966 228318 362146 228406
rect 362254 228318 362434 228406
rect 362542 228318 362722 228406
rect 362830 228318 363010 228406
rect 363264 228318 363444 228406
rect 363552 228318 363732 228406
rect 363840 228318 364020 228406
rect 364128 228318 364308 228406
rect 364416 228318 364596 228406
rect 364704 228318 364884 228406
rect 364992 228318 365172 228406
rect 365280 228318 365460 228406
rect 365714 228318 365894 228406
rect 366002 228318 366182 228406
rect 366290 228318 366470 228406
rect 366578 228318 366758 228406
rect 366866 228318 367046 228406
rect 367154 228318 367334 228406
rect 367442 228318 367622 228406
rect 367730 228318 367910 228406
rect 243214 228102 243394 228190
rect 243502 228102 243682 228190
rect 243790 228102 243970 228190
rect 244078 228102 244258 228190
rect 244366 228102 244546 228190
rect 244654 228102 244834 228190
rect 244942 228102 245122 228190
rect 245230 228102 245410 228190
rect 245664 228102 245844 228190
rect 245952 228102 246132 228190
rect 246240 228102 246420 228190
rect 246528 228102 246708 228190
rect 246816 228102 246996 228190
rect 247104 228102 247284 228190
rect 247392 228102 247572 228190
rect 247680 228102 247860 228190
rect 248114 228102 248294 228190
rect 248402 228102 248582 228190
rect 248690 228102 248870 228190
rect 248978 228102 249158 228190
rect 249266 228102 249446 228190
rect 249554 228102 249734 228190
rect 249842 228102 250022 228190
rect 250130 228102 250310 228190
rect 250564 228102 250744 228190
rect 360436 228102 360560 228190
rect 360814 228102 360994 228190
rect 361102 228102 361282 228190
rect 361390 228102 361570 228190
rect 361678 228102 361858 228190
rect 361966 228102 362146 228190
rect 362254 228102 362434 228190
rect 362542 228102 362722 228190
rect 362830 228102 363010 228190
rect 363264 228102 363444 228190
rect 363552 228102 363732 228190
rect 363840 228102 364020 228190
rect 364128 228102 364308 228190
rect 364416 228102 364596 228190
rect 364704 228102 364884 228190
rect 364992 228102 365172 228190
rect 365280 228102 365460 228190
rect 365714 228102 365894 228190
rect 366002 228102 366182 228190
rect 366290 228102 366470 228190
rect 366578 228102 366758 228190
rect 366866 228102 367046 228190
rect 367154 228102 367334 228190
rect 367442 228102 367622 228190
rect 367730 228102 367910 228190
rect 243214 227626 243394 227714
rect 243502 227626 243682 227714
rect 243790 227626 243970 227714
rect 244078 227626 244258 227714
rect 244366 227626 244546 227714
rect 244654 227626 244834 227714
rect 244942 227626 245122 227714
rect 245230 227626 245410 227714
rect 245664 227626 245844 227714
rect 245952 227626 246132 227714
rect 246240 227626 246420 227714
rect 246528 227626 246708 227714
rect 246816 227626 246996 227714
rect 247104 227626 247284 227714
rect 247392 227626 247572 227714
rect 247680 227626 247860 227714
rect 248114 227626 248294 227714
rect 248402 227626 248582 227714
rect 248690 227626 248870 227714
rect 248978 227626 249158 227714
rect 249266 227626 249446 227714
rect 249554 227626 249734 227714
rect 249842 227626 250022 227714
rect 250130 227626 250310 227714
rect 250564 227626 250744 227714
rect 360436 227626 360560 227714
rect 360814 227626 360994 227714
rect 361102 227626 361282 227714
rect 361390 227626 361570 227714
rect 361678 227626 361858 227714
rect 361966 227626 362146 227714
rect 362254 227626 362434 227714
rect 362542 227626 362722 227714
rect 362830 227626 363010 227714
rect 363264 227626 363444 227714
rect 363552 227626 363732 227714
rect 363840 227626 364020 227714
rect 364128 227626 364308 227714
rect 364416 227626 364596 227714
rect 364704 227626 364884 227714
rect 364992 227626 365172 227714
rect 365280 227626 365460 227714
rect 365714 227626 365894 227714
rect 366002 227626 366182 227714
rect 366290 227626 366470 227714
rect 366578 227626 366758 227714
rect 366866 227626 367046 227714
rect 367154 227626 367334 227714
rect 367442 227626 367622 227714
rect 367730 227626 367910 227714
rect 243214 227152 243394 227240
rect 243502 227152 243682 227240
rect 243790 227152 243970 227240
rect 244078 227152 244258 227240
rect 244366 227152 244546 227240
rect 244654 227152 244834 227240
rect 244942 227152 245122 227240
rect 245230 227152 245410 227240
rect 245664 227152 245844 227240
rect 245952 227152 246132 227240
rect 246240 227152 246420 227240
rect 246528 227152 246708 227240
rect 246816 227152 246996 227240
rect 247104 227152 247284 227240
rect 247392 227152 247572 227240
rect 247680 227152 247860 227240
rect 248114 227152 248294 227240
rect 248402 227152 248582 227240
rect 248690 227152 248870 227240
rect 248978 227152 249158 227240
rect 249266 227152 249446 227240
rect 249554 227152 249734 227240
rect 249842 227152 250022 227240
rect 250130 227152 250310 227240
rect 250564 227152 250744 227240
rect 360436 227152 360560 227240
rect 360814 227152 360994 227240
rect 361102 227152 361282 227240
rect 361390 227152 361570 227240
rect 361678 227152 361858 227240
rect 361966 227152 362146 227240
rect 362254 227152 362434 227240
rect 362542 227152 362722 227240
rect 362830 227152 363010 227240
rect 363264 227152 363444 227240
rect 363552 227152 363732 227240
rect 363840 227152 364020 227240
rect 364128 227152 364308 227240
rect 364416 227152 364596 227240
rect 364704 227152 364884 227240
rect 364992 227152 365172 227240
rect 365280 227152 365460 227240
rect 365714 227152 365894 227240
rect 366002 227152 366182 227240
rect 366290 227152 366470 227240
rect 366578 227152 366758 227240
rect 366866 227152 367046 227240
rect 367154 227152 367334 227240
rect 367442 227152 367622 227240
rect 367730 227152 367910 227240
rect 243214 226676 243394 226764
rect 243502 226676 243682 226764
rect 243790 226676 243970 226764
rect 244078 226676 244258 226764
rect 244366 226676 244546 226764
rect 244654 226676 244834 226764
rect 244942 226676 245122 226764
rect 245230 226676 245410 226764
rect 245664 226676 245844 226764
rect 245952 226676 246132 226764
rect 246240 226676 246420 226764
rect 246528 226676 246708 226764
rect 246816 226676 246996 226764
rect 247104 226676 247284 226764
rect 247392 226676 247572 226764
rect 247680 226676 247860 226764
rect 248114 226676 248294 226764
rect 248402 226676 248582 226764
rect 248690 226676 248870 226764
rect 248978 226676 249158 226764
rect 249266 226676 249446 226764
rect 249554 226676 249734 226764
rect 249842 226676 250022 226764
rect 250130 226676 250310 226764
rect 250564 226676 250744 226764
rect 360436 226676 360560 226764
rect 360814 226676 360994 226764
rect 361102 226676 361282 226764
rect 361390 226676 361570 226764
rect 361678 226676 361858 226764
rect 361966 226676 362146 226764
rect 362254 226676 362434 226764
rect 362542 226676 362722 226764
rect 362830 226676 363010 226764
rect 363264 226676 363444 226764
rect 363552 226676 363732 226764
rect 363840 226676 364020 226764
rect 364128 226676 364308 226764
rect 364416 226676 364596 226764
rect 364704 226676 364884 226764
rect 364992 226676 365172 226764
rect 365280 226676 365460 226764
rect 365714 226676 365894 226764
rect 366002 226676 366182 226764
rect 366290 226676 366470 226764
rect 366578 226676 366758 226764
rect 366866 226676 367046 226764
rect 367154 226676 367334 226764
rect 367442 226676 367622 226764
rect 367730 226676 367910 226764
rect 243214 226460 243394 226548
rect 243502 226460 243682 226548
rect 243790 226460 243970 226548
rect 244078 226460 244258 226548
rect 244366 226460 244546 226548
rect 244654 226460 244834 226548
rect 244942 226460 245122 226548
rect 245230 226460 245410 226548
rect 245664 226460 245844 226548
rect 245952 226460 246132 226548
rect 246240 226460 246420 226548
rect 246528 226460 246708 226548
rect 246816 226460 246996 226548
rect 247104 226460 247284 226548
rect 247392 226460 247572 226548
rect 247680 226460 247860 226548
rect 248114 226460 248294 226548
rect 248402 226460 248582 226548
rect 248690 226460 248870 226548
rect 248978 226460 249158 226548
rect 249266 226460 249446 226548
rect 249554 226460 249734 226548
rect 249842 226460 250022 226548
rect 250130 226460 250310 226548
rect 250564 226460 250744 226548
rect 360436 226460 360560 226548
rect 360814 226460 360994 226548
rect 361102 226460 361282 226548
rect 361390 226460 361570 226548
rect 361678 226460 361858 226548
rect 361966 226460 362146 226548
rect 362254 226460 362434 226548
rect 362542 226460 362722 226548
rect 362830 226460 363010 226548
rect 363264 226460 363444 226548
rect 363552 226460 363732 226548
rect 363840 226460 364020 226548
rect 364128 226460 364308 226548
rect 364416 226460 364596 226548
rect 364704 226460 364884 226548
rect 364992 226460 365172 226548
rect 365280 226460 365460 226548
rect 365714 226460 365894 226548
rect 366002 226460 366182 226548
rect 366290 226460 366470 226548
rect 366578 226460 366758 226548
rect 366866 226460 367046 226548
rect 367154 226460 367334 226548
rect 367442 226460 367622 226548
rect 367730 226460 367910 226548
rect 243214 225984 243394 226072
rect 243502 225984 243682 226072
rect 243790 225984 243970 226072
rect 244078 225984 244258 226072
rect 244366 225984 244546 226072
rect 244654 225984 244834 226072
rect 244942 225984 245122 226072
rect 245230 225984 245410 226072
rect 245664 225984 245844 226072
rect 245952 225984 246132 226072
rect 246240 225984 246420 226072
rect 246528 225984 246708 226072
rect 246816 225984 246996 226072
rect 247104 225984 247284 226072
rect 247392 225984 247572 226072
rect 247680 225984 247860 226072
rect 248114 225984 248294 226072
rect 248402 225984 248582 226072
rect 248690 225984 248870 226072
rect 248978 225984 249158 226072
rect 249266 225984 249446 226072
rect 249554 225984 249734 226072
rect 249842 225984 250022 226072
rect 250130 225984 250310 226072
rect 250564 225984 250744 226072
rect 360436 225984 360560 226072
rect 360814 225984 360994 226072
rect 361102 225984 361282 226072
rect 361390 225984 361570 226072
rect 361678 225984 361858 226072
rect 361966 225984 362146 226072
rect 362254 225984 362434 226072
rect 362542 225984 362722 226072
rect 362830 225984 363010 226072
rect 363264 225984 363444 226072
rect 363552 225984 363732 226072
rect 363840 225984 364020 226072
rect 364128 225984 364308 226072
rect 364416 225984 364596 226072
rect 364704 225984 364884 226072
rect 364992 225984 365172 226072
rect 365280 225984 365460 226072
rect 365714 225984 365894 226072
rect 366002 225984 366182 226072
rect 366290 225984 366470 226072
rect 366578 225984 366758 226072
rect 366866 225984 367046 226072
rect 367154 225984 367334 226072
rect 367442 225984 367622 226072
rect 367730 225984 367910 226072
rect 243214 225768 243394 225856
rect 243502 225768 243682 225856
rect 243790 225768 243970 225856
rect 244078 225768 244258 225856
rect 244366 225768 244546 225856
rect 244654 225768 244834 225856
rect 244942 225768 245122 225856
rect 245230 225768 245410 225856
rect 245664 225768 245844 225856
rect 245952 225768 246132 225856
rect 246240 225768 246420 225856
rect 246528 225768 246708 225856
rect 246816 225768 246996 225856
rect 247104 225768 247284 225856
rect 247392 225768 247572 225856
rect 247680 225768 247860 225856
rect 248114 225768 248294 225856
rect 248402 225768 248582 225856
rect 248690 225768 248870 225856
rect 248978 225768 249158 225856
rect 249266 225768 249446 225856
rect 249554 225768 249734 225856
rect 249842 225768 250022 225856
rect 250130 225768 250310 225856
rect 250564 225768 250744 225856
rect 360436 225768 360560 225856
rect 360814 225768 360994 225856
rect 361102 225768 361282 225856
rect 361390 225768 361570 225856
rect 361678 225768 361858 225856
rect 361966 225768 362146 225856
rect 362254 225768 362434 225856
rect 362542 225768 362722 225856
rect 362830 225768 363010 225856
rect 363264 225768 363444 225856
rect 363552 225768 363732 225856
rect 363840 225768 364020 225856
rect 364128 225768 364308 225856
rect 364416 225768 364596 225856
rect 364704 225768 364884 225856
rect 364992 225768 365172 225856
rect 365280 225768 365460 225856
rect 365714 225768 365894 225856
rect 366002 225768 366182 225856
rect 366290 225768 366470 225856
rect 366578 225768 366758 225856
rect 366866 225768 367046 225856
rect 367154 225768 367334 225856
rect 367442 225768 367622 225856
rect 367730 225768 367910 225856
rect 243214 225292 243394 225380
rect 243502 225292 243682 225380
rect 243790 225292 243970 225380
rect 244078 225292 244258 225380
rect 244366 225292 244546 225380
rect 244654 225292 244834 225380
rect 244942 225292 245122 225380
rect 245230 225292 245410 225380
rect 245664 225292 245844 225380
rect 245952 225292 246132 225380
rect 246240 225292 246420 225380
rect 246528 225292 246708 225380
rect 246816 225292 246996 225380
rect 247104 225292 247284 225380
rect 247392 225292 247572 225380
rect 247680 225292 247860 225380
rect 248114 225292 248294 225380
rect 248402 225292 248582 225380
rect 248690 225292 248870 225380
rect 248978 225292 249158 225380
rect 249266 225292 249446 225380
rect 249554 225292 249734 225380
rect 249842 225292 250022 225380
rect 250130 225292 250310 225380
rect 250564 225292 250744 225380
rect 360436 225292 360560 225380
rect 360814 225292 360994 225380
rect 361102 225292 361282 225380
rect 361390 225292 361570 225380
rect 361678 225292 361858 225380
rect 361966 225292 362146 225380
rect 362254 225292 362434 225380
rect 362542 225292 362722 225380
rect 362830 225292 363010 225380
rect 363264 225292 363444 225380
rect 363552 225292 363732 225380
rect 363840 225292 364020 225380
rect 364128 225292 364308 225380
rect 364416 225292 364596 225380
rect 364704 225292 364884 225380
rect 364992 225292 365172 225380
rect 365280 225292 365460 225380
rect 365714 225292 365894 225380
rect 366002 225292 366182 225380
rect 366290 225292 366470 225380
rect 366578 225292 366758 225380
rect 366866 225292 367046 225380
rect 367154 225292 367334 225380
rect 367442 225292 367622 225380
rect 367730 225292 367910 225380
rect 243214 225076 243394 225164
rect 243502 225076 243682 225164
rect 243790 225076 243970 225164
rect 244078 225076 244258 225164
rect 244366 225076 244546 225164
rect 244654 225076 244834 225164
rect 244942 225076 245122 225164
rect 245230 225076 245410 225164
rect 245664 225076 245844 225164
rect 245952 225076 246132 225164
rect 246240 225076 246420 225164
rect 246528 225076 246708 225164
rect 246816 225076 246996 225164
rect 247104 225076 247284 225164
rect 247392 225076 247572 225164
rect 247680 225076 247860 225164
rect 248114 225076 248294 225164
rect 248402 225076 248582 225164
rect 248690 225076 248870 225164
rect 248978 225076 249158 225164
rect 249266 225076 249446 225164
rect 249554 225076 249734 225164
rect 249842 225076 250022 225164
rect 250130 225076 250310 225164
rect 250564 225076 250744 225164
rect 360436 225076 360560 225164
rect 360814 225076 360994 225164
rect 361102 225076 361282 225164
rect 361390 225076 361570 225164
rect 361678 225076 361858 225164
rect 361966 225076 362146 225164
rect 362254 225076 362434 225164
rect 362542 225076 362722 225164
rect 362830 225076 363010 225164
rect 363264 225076 363444 225164
rect 363552 225076 363732 225164
rect 363840 225076 364020 225164
rect 364128 225076 364308 225164
rect 364416 225076 364596 225164
rect 364704 225076 364884 225164
rect 364992 225076 365172 225164
rect 365280 225076 365460 225164
rect 365714 225076 365894 225164
rect 366002 225076 366182 225164
rect 366290 225076 366470 225164
rect 366578 225076 366758 225164
rect 366866 225076 367046 225164
rect 367154 225076 367334 225164
rect 367442 225076 367622 225164
rect 367730 225076 367910 225164
rect 243214 224600 243394 224688
rect 243502 224600 243682 224688
rect 243790 224600 243970 224688
rect 244078 224600 244258 224688
rect 244366 224600 244546 224688
rect 244654 224600 244834 224688
rect 244942 224600 245122 224688
rect 245230 224600 245410 224688
rect 245664 224600 245844 224688
rect 245952 224600 246132 224688
rect 246240 224600 246420 224688
rect 246528 224600 246708 224688
rect 246816 224600 246996 224688
rect 247104 224600 247284 224688
rect 247392 224600 247572 224688
rect 247680 224600 247860 224688
rect 248114 224600 248294 224688
rect 248402 224600 248582 224688
rect 248690 224600 248870 224688
rect 248978 224600 249158 224688
rect 249266 224600 249446 224688
rect 249554 224600 249734 224688
rect 249842 224600 250022 224688
rect 250130 224600 250310 224688
rect 250564 224600 250744 224688
rect 360436 224600 360560 224688
rect 360814 224600 360994 224688
rect 361102 224600 361282 224688
rect 361390 224600 361570 224688
rect 361678 224600 361858 224688
rect 361966 224600 362146 224688
rect 362254 224600 362434 224688
rect 362542 224600 362722 224688
rect 362830 224600 363010 224688
rect 363264 224600 363444 224688
rect 363552 224600 363732 224688
rect 363840 224600 364020 224688
rect 364128 224600 364308 224688
rect 364416 224600 364596 224688
rect 364704 224600 364884 224688
rect 364992 224600 365172 224688
rect 365280 224600 365460 224688
rect 365714 224600 365894 224688
rect 366002 224600 366182 224688
rect 366290 224600 366470 224688
rect 366578 224600 366758 224688
rect 366866 224600 367046 224688
rect 367154 224600 367334 224688
rect 367442 224600 367622 224688
rect 367730 224600 367910 224688
rect 243214 224126 243394 224214
rect 243502 224126 243682 224214
rect 243790 224126 243970 224214
rect 244078 224126 244258 224214
rect 244366 224126 244546 224214
rect 244654 224126 244834 224214
rect 244942 224126 245122 224214
rect 245230 224126 245410 224214
rect 245664 224126 245844 224214
rect 245952 224126 246132 224214
rect 246240 224126 246420 224214
rect 246528 224126 246708 224214
rect 246816 224126 246996 224214
rect 247104 224126 247284 224214
rect 247392 224126 247572 224214
rect 247680 224126 247860 224214
rect 248114 224126 248294 224214
rect 248402 224126 248582 224214
rect 248690 224126 248870 224214
rect 248978 224126 249158 224214
rect 249266 224126 249446 224214
rect 249554 224126 249734 224214
rect 249842 224126 250022 224214
rect 250130 224126 250310 224214
rect 250564 224126 250744 224214
rect 360436 224126 360560 224214
rect 360814 224126 360994 224214
rect 361102 224126 361282 224214
rect 361390 224126 361570 224214
rect 361678 224126 361858 224214
rect 361966 224126 362146 224214
rect 362254 224126 362434 224214
rect 362542 224126 362722 224214
rect 362830 224126 363010 224214
rect 363264 224126 363444 224214
rect 363552 224126 363732 224214
rect 363840 224126 364020 224214
rect 364128 224126 364308 224214
rect 364416 224126 364596 224214
rect 364704 224126 364884 224214
rect 364992 224126 365172 224214
rect 365280 224126 365460 224214
rect 365714 224126 365894 224214
rect 366002 224126 366182 224214
rect 366290 224126 366470 224214
rect 366578 224126 366758 224214
rect 366866 224126 367046 224214
rect 367154 224126 367334 224214
rect 367442 224126 367622 224214
rect 367730 224126 367910 224214
rect 243214 223650 243394 223738
rect 243502 223650 243682 223738
rect 243790 223650 243970 223738
rect 244078 223650 244258 223738
rect 244366 223650 244546 223738
rect 244654 223650 244834 223738
rect 244942 223650 245122 223738
rect 245230 223650 245410 223738
rect 245664 223650 245844 223738
rect 245952 223650 246132 223738
rect 246240 223650 246420 223738
rect 246528 223650 246708 223738
rect 246816 223650 246996 223738
rect 247104 223650 247284 223738
rect 247392 223650 247572 223738
rect 247680 223650 247860 223738
rect 248114 223650 248294 223738
rect 248402 223650 248582 223738
rect 248690 223650 248870 223738
rect 248978 223650 249158 223738
rect 249266 223650 249446 223738
rect 249554 223650 249734 223738
rect 249842 223650 250022 223738
rect 250130 223650 250310 223738
rect 250564 223650 250744 223738
rect 360436 223650 360560 223738
rect 360814 223650 360994 223738
rect 361102 223650 361282 223738
rect 361390 223650 361570 223738
rect 361678 223650 361858 223738
rect 361966 223650 362146 223738
rect 362254 223650 362434 223738
rect 362542 223650 362722 223738
rect 362830 223650 363010 223738
rect 363264 223650 363444 223738
rect 363552 223650 363732 223738
rect 363840 223650 364020 223738
rect 364128 223650 364308 223738
rect 364416 223650 364596 223738
rect 364704 223650 364884 223738
rect 364992 223650 365172 223738
rect 365280 223650 365460 223738
rect 365714 223650 365894 223738
rect 366002 223650 366182 223738
rect 366290 223650 366470 223738
rect 366578 223650 366758 223738
rect 366866 223650 367046 223738
rect 367154 223650 367334 223738
rect 367442 223650 367622 223738
rect 367730 223650 367910 223738
rect 243214 223434 243394 223522
rect 243502 223434 243682 223522
rect 243790 223434 243970 223522
rect 244078 223434 244258 223522
rect 244366 223434 244546 223522
rect 244654 223434 244834 223522
rect 244942 223434 245122 223522
rect 245230 223434 245410 223522
rect 245664 223434 245844 223522
rect 245952 223434 246132 223522
rect 246240 223434 246420 223522
rect 246528 223434 246708 223522
rect 246816 223434 246996 223522
rect 247104 223434 247284 223522
rect 247392 223434 247572 223522
rect 247680 223434 247860 223522
rect 248114 223434 248294 223522
rect 248402 223434 248582 223522
rect 248690 223434 248870 223522
rect 248978 223434 249158 223522
rect 249266 223434 249446 223522
rect 249554 223434 249734 223522
rect 249842 223434 250022 223522
rect 250130 223434 250310 223522
rect 250564 223434 250744 223522
rect 360436 223434 360560 223522
rect 360814 223434 360994 223522
rect 361102 223434 361282 223522
rect 361390 223434 361570 223522
rect 361678 223434 361858 223522
rect 361966 223434 362146 223522
rect 362254 223434 362434 223522
rect 362542 223434 362722 223522
rect 362830 223434 363010 223522
rect 363264 223434 363444 223522
rect 363552 223434 363732 223522
rect 363840 223434 364020 223522
rect 364128 223434 364308 223522
rect 364416 223434 364596 223522
rect 364704 223434 364884 223522
rect 364992 223434 365172 223522
rect 365280 223434 365460 223522
rect 365714 223434 365894 223522
rect 366002 223434 366182 223522
rect 366290 223434 366470 223522
rect 366578 223434 366758 223522
rect 366866 223434 367046 223522
rect 367154 223434 367334 223522
rect 367442 223434 367622 223522
rect 367730 223434 367910 223522
rect 243214 222958 243394 223046
rect 243502 222958 243682 223046
rect 243790 222958 243970 223046
rect 244078 222958 244258 223046
rect 244366 222958 244546 223046
rect 244654 222958 244834 223046
rect 244942 222958 245122 223046
rect 245230 222958 245410 223046
rect 245664 222958 245844 223046
rect 245952 222958 246132 223046
rect 246240 222958 246420 223046
rect 246528 222958 246708 223046
rect 246816 222958 246996 223046
rect 247104 222958 247284 223046
rect 247392 222958 247572 223046
rect 247680 222958 247860 223046
rect 248114 222958 248294 223046
rect 248402 222958 248582 223046
rect 248690 222958 248870 223046
rect 248978 222958 249158 223046
rect 249266 222958 249446 223046
rect 249554 222958 249734 223046
rect 249842 222958 250022 223046
rect 250130 222958 250310 223046
rect 250564 222958 250744 223046
rect 360436 222958 360560 223046
rect 360814 222958 360994 223046
rect 361102 222958 361282 223046
rect 361390 222958 361570 223046
rect 361678 222958 361858 223046
rect 361966 222958 362146 223046
rect 362254 222958 362434 223046
rect 362542 222958 362722 223046
rect 362830 222958 363010 223046
rect 363264 222958 363444 223046
rect 363552 222958 363732 223046
rect 363840 222958 364020 223046
rect 364128 222958 364308 223046
rect 364416 222958 364596 223046
rect 364704 222958 364884 223046
rect 364992 222958 365172 223046
rect 365280 222958 365460 223046
rect 365714 222958 365894 223046
rect 366002 222958 366182 223046
rect 366290 222958 366470 223046
rect 366578 222958 366758 223046
rect 366866 222958 367046 223046
rect 367154 222958 367334 223046
rect 367442 222958 367622 223046
rect 367730 222958 367910 223046
rect 243214 222742 243394 222830
rect 243502 222742 243682 222830
rect 243790 222742 243970 222830
rect 244078 222742 244258 222830
rect 244366 222742 244546 222830
rect 244654 222742 244834 222830
rect 244942 222742 245122 222830
rect 245230 222742 245410 222830
rect 245664 222742 245844 222830
rect 245952 222742 246132 222830
rect 246240 222742 246420 222830
rect 246528 222742 246708 222830
rect 246816 222742 246996 222830
rect 247104 222742 247284 222830
rect 247392 222742 247572 222830
rect 247680 222742 247860 222830
rect 248114 222742 248294 222830
rect 248402 222742 248582 222830
rect 248690 222742 248870 222830
rect 248978 222742 249158 222830
rect 249266 222742 249446 222830
rect 249554 222742 249734 222830
rect 249842 222742 250022 222830
rect 250130 222742 250310 222830
rect 250564 222742 250744 222830
rect 360436 222742 360560 222830
rect 360814 222742 360994 222830
rect 361102 222742 361282 222830
rect 361390 222742 361570 222830
rect 361678 222742 361858 222830
rect 361966 222742 362146 222830
rect 362254 222742 362434 222830
rect 362542 222742 362722 222830
rect 362830 222742 363010 222830
rect 363264 222742 363444 222830
rect 363552 222742 363732 222830
rect 363840 222742 364020 222830
rect 364128 222742 364308 222830
rect 364416 222742 364596 222830
rect 364704 222742 364884 222830
rect 364992 222742 365172 222830
rect 365280 222742 365460 222830
rect 365714 222742 365894 222830
rect 366002 222742 366182 222830
rect 366290 222742 366470 222830
rect 366578 222742 366758 222830
rect 366866 222742 367046 222830
rect 367154 222742 367334 222830
rect 367442 222742 367622 222830
rect 367730 222742 367910 222830
rect 243214 222266 243394 222354
rect 243502 222266 243682 222354
rect 243790 222266 243970 222354
rect 244078 222266 244258 222354
rect 244366 222266 244546 222354
rect 244654 222266 244834 222354
rect 244942 222266 245122 222354
rect 245230 222266 245410 222354
rect 245664 222266 245844 222354
rect 245952 222266 246132 222354
rect 246240 222266 246420 222354
rect 246528 222266 246708 222354
rect 246816 222266 246996 222354
rect 247104 222266 247284 222354
rect 247392 222266 247572 222354
rect 247680 222266 247860 222354
rect 248114 222266 248294 222354
rect 248402 222266 248582 222354
rect 248690 222266 248870 222354
rect 248978 222266 249158 222354
rect 249266 222266 249446 222354
rect 249554 222266 249734 222354
rect 249842 222266 250022 222354
rect 250130 222266 250310 222354
rect 250564 222266 250744 222354
rect 360436 222266 360560 222354
rect 360814 222266 360994 222354
rect 361102 222266 361282 222354
rect 361390 222266 361570 222354
rect 361678 222266 361858 222354
rect 361966 222266 362146 222354
rect 362254 222266 362434 222354
rect 362542 222266 362722 222354
rect 362830 222266 363010 222354
rect 363264 222266 363444 222354
rect 363552 222266 363732 222354
rect 363840 222266 364020 222354
rect 364128 222266 364308 222354
rect 364416 222266 364596 222354
rect 364704 222266 364884 222354
rect 364992 222266 365172 222354
rect 365280 222266 365460 222354
rect 365714 222266 365894 222354
rect 366002 222266 366182 222354
rect 366290 222266 366470 222354
rect 366578 222266 366758 222354
rect 366866 222266 367046 222354
rect 367154 222266 367334 222354
rect 367442 222266 367622 222354
rect 367730 222266 367910 222354
rect 243214 222050 243394 222138
rect 243502 222050 243682 222138
rect 243790 222050 243970 222138
rect 244078 222050 244258 222138
rect 244366 222050 244546 222138
rect 244654 222050 244834 222138
rect 244942 222050 245122 222138
rect 245230 222050 245410 222138
rect 245664 222050 245844 222138
rect 245952 222050 246132 222138
rect 246240 222050 246420 222138
rect 246528 222050 246708 222138
rect 246816 222050 246996 222138
rect 247104 222050 247284 222138
rect 247392 222050 247572 222138
rect 247680 222050 247860 222138
rect 248114 222050 248294 222138
rect 248402 222050 248582 222138
rect 248690 222050 248870 222138
rect 248978 222050 249158 222138
rect 249266 222050 249446 222138
rect 249554 222050 249734 222138
rect 249842 222050 250022 222138
rect 250130 222050 250310 222138
rect 250564 222050 250744 222138
rect 360436 222050 360560 222138
rect 360814 222050 360994 222138
rect 361102 222050 361282 222138
rect 361390 222050 361570 222138
rect 361678 222050 361858 222138
rect 361966 222050 362146 222138
rect 362254 222050 362434 222138
rect 362542 222050 362722 222138
rect 362830 222050 363010 222138
rect 363264 222050 363444 222138
rect 363552 222050 363732 222138
rect 363840 222050 364020 222138
rect 364128 222050 364308 222138
rect 364416 222050 364596 222138
rect 364704 222050 364884 222138
rect 364992 222050 365172 222138
rect 365280 222050 365460 222138
rect 365714 222050 365894 222138
rect 366002 222050 366182 222138
rect 366290 222050 366470 222138
rect 366578 222050 366758 222138
rect 366866 222050 367046 222138
rect 367154 222050 367334 222138
rect 367442 222050 367622 222138
rect 367730 222050 367910 222138
rect 243214 221574 243394 221662
rect 243502 221574 243682 221662
rect 243790 221574 243970 221662
rect 244078 221574 244258 221662
rect 244366 221574 244546 221662
rect 244654 221574 244834 221662
rect 244942 221574 245122 221662
rect 245230 221574 245410 221662
rect 245664 221574 245844 221662
rect 245952 221574 246132 221662
rect 246240 221574 246420 221662
rect 246528 221574 246708 221662
rect 246816 221574 246996 221662
rect 247104 221574 247284 221662
rect 247392 221574 247572 221662
rect 247680 221574 247860 221662
rect 248114 221574 248294 221662
rect 248402 221574 248582 221662
rect 248690 221574 248870 221662
rect 248978 221574 249158 221662
rect 249266 221574 249446 221662
rect 249554 221574 249734 221662
rect 249842 221574 250022 221662
rect 250130 221574 250310 221662
rect 250564 221574 250744 221662
rect 360436 221574 360560 221662
rect 360814 221574 360994 221662
rect 361102 221574 361282 221662
rect 361390 221574 361570 221662
rect 361678 221574 361858 221662
rect 361966 221574 362146 221662
rect 362254 221574 362434 221662
rect 362542 221574 362722 221662
rect 362830 221574 363010 221662
rect 363264 221574 363444 221662
rect 363552 221574 363732 221662
rect 363840 221574 364020 221662
rect 364128 221574 364308 221662
rect 364416 221574 364596 221662
rect 364704 221574 364884 221662
rect 364992 221574 365172 221662
rect 365280 221574 365460 221662
rect 365714 221574 365894 221662
rect 366002 221574 366182 221662
rect 366290 221574 366470 221662
rect 366578 221574 366758 221662
rect 366866 221574 367046 221662
rect 367154 221574 367334 221662
rect 367442 221574 367622 221662
rect 367730 221574 367910 221662
rect 243214 221100 243394 221188
rect 243502 221100 243682 221188
rect 243790 221100 243970 221188
rect 244078 221100 244258 221188
rect 244366 221100 244546 221188
rect 244654 221100 244834 221188
rect 244942 221100 245122 221188
rect 245230 221100 245410 221188
rect 245664 221100 245844 221188
rect 245952 221100 246132 221188
rect 246240 221100 246420 221188
rect 246528 221100 246708 221188
rect 246816 221100 246996 221188
rect 247104 221100 247284 221188
rect 247392 221100 247572 221188
rect 247680 221100 247860 221188
rect 248114 221100 248294 221188
rect 248402 221100 248582 221188
rect 248690 221100 248870 221188
rect 248978 221100 249158 221188
rect 249266 221100 249446 221188
rect 249554 221100 249734 221188
rect 249842 221100 250022 221188
rect 250130 221100 250310 221188
rect 250564 221100 250744 221188
rect 360436 221100 360560 221188
rect 360814 221100 360994 221188
rect 361102 221100 361282 221188
rect 361390 221100 361570 221188
rect 361678 221100 361858 221188
rect 361966 221100 362146 221188
rect 362254 221100 362434 221188
rect 362542 221100 362722 221188
rect 362830 221100 363010 221188
rect 363264 221100 363444 221188
rect 363552 221100 363732 221188
rect 363840 221100 364020 221188
rect 364128 221100 364308 221188
rect 364416 221100 364596 221188
rect 364704 221100 364884 221188
rect 364992 221100 365172 221188
rect 365280 221100 365460 221188
rect 365714 221100 365894 221188
rect 366002 221100 366182 221188
rect 366290 221100 366470 221188
rect 366578 221100 366758 221188
rect 366866 221100 367046 221188
rect 367154 221100 367334 221188
rect 367442 221100 367622 221188
rect 367730 221100 367910 221188
rect 243214 220624 243394 220712
rect 243502 220624 243682 220712
rect 243790 220624 243970 220712
rect 244078 220624 244258 220712
rect 244366 220624 244546 220712
rect 244654 220624 244834 220712
rect 244942 220624 245122 220712
rect 245230 220624 245410 220712
rect 245664 220624 245844 220712
rect 245952 220624 246132 220712
rect 246240 220624 246420 220712
rect 246528 220624 246708 220712
rect 246816 220624 246996 220712
rect 247104 220624 247284 220712
rect 247392 220624 247572 220712
rect 247680 220624 247860 220712
rect 248114 220624 248294 220712
rect 248402 220624 248582 220712
rect 248690 220624 248870 220712
rect 248978 220624 249158 220712
rect 249266 220624 249446 220712
rect 249554 220624 249734 220712
rect 249842 220624 250022 220712
rect 250130 220624 250310 220712
rect 250564 220624 250744 220712
rect 360436 220624 360560 220712
rect 360814 220624 360994 220712
rect 361102 220624 361282 220712
rect 361390 220624 361570 220712
rect 361678 220624 361858 220712
rect 361966 220624 362146 220712
rect 362254 220624 362434 220712
rect 362542 220624 362722 220712
rect 362830 220624 363010 220712
rect 363264 220624 363444 220712
rect 363552 220624 363732 220712
rect 363840 220624 364020 220712
rect 364128 220624 364308 220712
rect 364416 220624 364596 220712
rect 364704 220624 364884 220712
rect 364992 220624 365172 220712
rect 365280 220624 365460 220712
rect 365714 220624 365894 220712
rect 366002 220624 366182 220712
rect 366290 220624 366470 220712
rect 366578 220624 366758 220712
rect 366866 220624 367046 220712
rect 367154 220624 367334 220712
rect 367442 220624 367622 220712
rect 367730 220624 367910 220712
rect 243214 220408 243394 220496
rect 243502 220408 243682 220496
rect 243790 220408 243970 220496
rect 244078 220408 244258 220496
rect 244366 220408 244546 220496
rect 244654 220408 244834 220496
rect 244942 220408 245122 220496
rect 245230 220408 245410 220496
rect 245664 220408 245844 220496
rect 245952 220408 246132 220496
rect 246240 220408 246420 220496
rect 246528 220408 246708 220496
rect 246816 220408 246996 220496
rect 247104 220408 247284 220496
rect 247392 220408 247572 220496
rect 247680 220408 247860 220496
rect 248114 220408 248294 220496
rect 248402 220408 248582 220496
rect 248690 220408 248870 220496
rect 248978 220408 249158 220496
rect 249266 220408 249446 220496
rect 249554 220408 249734 220496
rect 249842 220408 250022 220496
rect 250130 220408 250310 220496
rect 250564 220408 250744 220496
rect 360436 220408 360560 220496
rect 360814 220408 360994 220496
rect 361102 220408 361282 220496
rect 361390 220408 361570 220496
rect 361678 220408 361858 220496
rect 361966 220408 362146 220496
rect 362254 220408 362434 220496
rect 362542 220408 362722 220496
rect 362830 220408 363010 220496
rect 363264 220408 363444 220496
rect 363552 220408 363732 220496
rect 363840 220408 364020 220496
rect 364128 220408 364308 220496
rect 364416 220408 364596 220496
rect 364704 220408 364884 220496
rect 364992 220408 365172 220496
rect 365280 220408 365460 220496
rect 365714 220408 365894 220496
rect 366002 220408 366182 220496
rect 366290 220408 366470 220496
rect 366578 220408 366758 220496
rect 366866 220408 367046 220496
rect 367154 220408 367334 220496
rect 367442 220408 367622 220496
rect 367730 220408 367910 220496
rect 243214 219932 243394 220020
rect 243502 219932 243682 220020
rect 243790 219932 243970 220020
rect 244078 219932 244258 220020
rect 244366 219932 244546 220020
rect 244654 219932 244834 220020
rect 244942 219932 245122 220020
rect 245230 219932 245410 220020
rect 245664 219932 245844 220020
rect 245952 219932 246132 220020
rect 246240 219932 246420 220020
rect 246528 219932 246708 220020
rect 246816 219932 246996 220020
rect 247104 219932 247284 220020
rect 247392 219932 247572 220020
rect 247680 219932 247860 220020
rect 248114 219932 248294 220020
rect 248402 219932 248582 220020
rect 248690 219932 248870 220020
rect 248978 219932 249158 220020
rect 249266 219932 249446 220020
rect 249554 219932 249734 220020
rect 249842 219932 250022 220020
rect 250130 219932 250310 220020
rect 250564 219932 250744 220020
rect 360436 219932 360560 220020
rect 360814 219932 360994 220020
rect 361102 219932 361282 220020
rect 361390 219932 361570 220020
rect 361678 219932 361858 220020
rect 361966 219932 362146 220020
rect 362254 219932 362434 220020
rect 362542 219932 362722 220020
rect 362830 219932 363010 220020
rect 363264 219932 363444 220020
rect 363552 219932 363732 220020
rect 363840 219932 364020 220020
rect 364128 219932 364308 220020
rect 364416 219932 364596 220020
rect 364704 219932 364884 220020
rect 364992 219932 365172 220020
rect 365280 219932 365460 220020
rect 365714 219932 365894 220020
rect 366002 219932 366182 220020
rect 366290 219932 366470 220020
rect 366578 219932 366758 220020
rect 366866 219932 367046 220020
rect 367154 219932 367334 220020
rect 367442 219932 367622 220020
rect 367730 219932 367910 220020
rect 243214 219716 243394 219804
rect 243502 219716 243682 219804
rect 243790 219716 243970 219804
rect 244078 219716 244258 219804
rect 244366 219716 244546 219804
rect 244654 219716 244834 219804
rect 244942 219716 245122 219804
rect 245230 219716 245410 219804
rect 245664 219716 245844 219804
rect 245952 219716 246132 219804
rect 246240 219716 246420 219804
rect 246528 219716 246708 219804
rect 246816 219716 246996 219804
rect 247104 219716 247284 219804
rect 247392 219716 247572 219804
rect 247680 219716 247860 219804
rect 248114 219716 248294 219804
rect 248402 219716 248582 219804
rect 248690 219716 248870 219804
rect 248978 219716 249158 219804
rect 249266 219716 249446 219804
rect 249554 219716 249734 219804
rect 249842 219716 250022 219804
rect 250130 219716 250310 219804
rect 250564 219716 250744 219804
rect 360436 219716 360560 219804
rect 360814 219716 360994 219804
rect 361102 219716 361282 219804
rect 361390 219716 361570 219804
rect 361678 219716 361858 219804
rect 361966 219716 362146 219804
rect 362254 219716 362434 219804
rect 362542 219716 362722 219804
rect 362830 219716 363010 219804
rect 363264 219716 363444 219804
rect 363552 219716 363732 219804
rect 363840 219716 364020 219804
rect 364128 219716 364308 219804
rect 364416 219716 364596 219804
rect 364704 219716 364884 219804
rect 364992 219716 365172 219804
rect 365280 219716 365460 219804
rect 365714 219716 365894 219804
rect 366002 219716 366182 219804
rect 366290 219716 366470 219804
rect 366578 219716 366758 219804
rect 366866 219716 367046 219804
rect 367154 219716 367334 219804
rect 367442 219716 367622 219804
rect 367730 219716 367910 219804
rect 243214 219240 243394 219328
rect 243502 219240 243682 219328
rect 243790 219240 243970 219328
rect 244078 219240 244258 219328
rect 244366 219240 244546 219328
rect 244654 219240 244834 219328
rect 244942 219240 245122 219328
rect 245230 219240 245410 219328
rect 245664 219240 245844 219328
rect 245952 219240 246132 219328
rect 246240 219240 246420 219328
rect 246528 219240 246708 219328
rect 246816 219240 246996 219328
rect 247104 219240 247284 219328
rect 247392 219240 247572 219328
rect 247680 219240 247860 219328
rect 248114 219240 248294 219328
rect 248402 219240 248582 219328
rect 248690 219240 248870 219328
rect 248978 219240 249158 219328
rect 249266 219240 249446 219328
rect 249554 219240 249734 219328
rect 249842 219240 250022 219328
rect 250130 219240 250310 219328
rect 250564 219240 250744 219328
rect 360436 219240 360560 219328
rect 360814 219240 360994 219328
rect 361102 219240 361282 219328
rect 361390 219240 361570 219328
rect 361678 219240 361858 219328
rect 361966 219240 362146 219328
rect 362254 219240 362434 219328
rect 362542 219240 362722 219328
rect 362830 219240 363010 219328
rect 363264 219240 363444 219328
rect 363552 219240 363732 219328
rect 363840 219240 364020 219328
rect 364128 219240 364308 219328
rect 364416 219240 364596 219328
rect 364704 219240 364884 219328
rect 364992 219240 365172 219328
rect 365280 219240 365460 219328
rect 365714 219240 365894 219328
rect 366002 219240 366182 219328
rect 366290 219240 366470 219328
rect 366578 219240 366758 219328
rect 366866 219240 367046 219328
rect 367154 219240 367334 219328
rect 367442 219240 367622 219328
rect 367730 219240 367910 219328
rect 243214 219024 243394 219112
rect 243502 219024 243682 219112
rect 243790 219024 243970 219112
rect 244078 219024 244258 219112
rect 244366 219024 244546 219112
rect 244654 219024 244834 219112
rect 244942 219024 245122 219112
rect 245230 219024 245410 219112
rect 245664 219024 245844 219112
rect 245952 219024 246132 219112
rect 246240 219024 246420 219112
rect 246528 219024 246708 219112
rect 246816 219024 246996 219112
rect 247104 219024 247284 219112
rect 247392 219024 247572 219112
rect 247680 219024 247860 219112
rect 248114 219024 248294 219112
rect 248402 219024 248582 219112
rect 248690 219024 248870 219112
rect 248978 219024 249158 219112
rect 249266 219024 249446 219112
rect 249554 219024 249734 219112
rect 249842 219024 250022 219112
rect 250130 219024 250310 219112
rect 250564 219024 250744 219112
rect 360436 219024 360560 219112
rect 360814 219024 360994 219112
rect 361102 219024 361282 219112
rect 361390 219024 361570 219112
rect 361678 219024 361858 219112
rect 361966 219024 362146 219112
rect 362254 219024 362434 219112
rect 362542 219024 362722 219112
rect 362830 219024 363010 219112
rect 363264 219024 363444 219112
rect 363552 219024 363732 219112
rect 363840 219024 364020 219112
rect 364128 219024 364308 219112
rect 364416 219024 364596 219112
rect 364704 219024 364884 219112
rect 364992 219024 365172 219112
rect 365280 219024 365460 219112
rect 365714 219024 365894 219112
rect 366002 219024 366182 219112
rect 366290 219024 366470 219112
rect 366578 219024 366758 219112
rect 366866 219024 367046 219112
rect 367154 219024 367334 219112
rect 367442 219024 367622 219112
rect 367730 219024 367910 219112
rect 243214 218548 243394 218636
rect 243502 218548 243682 218636
rect 243790 218548 243970 218636
rect 244078 218548 244258 218636
rect 244366 218548 244546 218636
rect 244654 218548 244834 218636
rect 244942 218548 245122 218636
rect 245230 218548 245410 218636
rect 245664 218548 245844 218636
rect 245952 218548 246132 218636
rect 246240 218548 246420 218636
rect 246528 218548 246708 218636
rect 246816 218548 246996 218636
rect 247104 218548 247284 218636
rect 247392 218548 247572 218636
rect 247680 218548 247860 218636
rect 248114 218548 248294 218636
rect 248402 218548 248582 218636
rect 248690 218548 248870 218636
rect 248978 218548 249158 218636
rect 249266 218548 249446 218636
rect 249554 218548 249734 218636
rect 249842 218548 250022 218636
rect 250130 218548 250310 218636
rect 250564 218548 250744 218636
rect 360436 218548 360560 218636
rect 360814 218548 360994 218636
rect 361102 218548 361282 218636
rect 361390 218548 361570 218636
rect 361678 218548 361858 218636
rect 361966 218548 362146 218636
rect 362254 218548 362434 218636
rect 362542 218548 362722 218636
rect 362830 218548 363010 218636
rect 363264 218548 363444 218636
rect 363552 218548 363732 218636
rect 363840 218548 364020 218636
rect 364128 218548 364308 218636
rect 364416 218548 364596 218636
rect 364704 218548 364884 218636
rect 364992 218548 365172 218636
rect 365280 218548 365460 218636
rect 365714 218548 365894 218636
rect 366002 218548 366182 218636
rect 366290 218548 366470 218636
rect 366578 218548 366758 218636
rect 366866 218548 367046 218636
rect 367154 218548 367334 218636
rect 367442 218548 367622 218636
rect 367730 218548 367910 218636
rect 243214 218074 243394 218162
rect 243502 218074 243682 218162
rect 243790 218074 243970 218162
rect 244078 218074 244258 218162
rect 244366 218074 244546 218162
rect 244654 218074 244834 218162
rect 244942 218074 245122 218162
rect 245230 218074 245410 218162
rect 245664 218074 245844 218162
rect 245952 218074 246132 218162
rect 246240 218074 246420 218162
rect 246528 218074 246708 218162
rect 246816 218074 246996 218162
rect 247104 218074 247284 218162
rect 247392 218074 247572 218162
rect 247680 218074 247860 218162
rect 248114 218074 248294 218162
rect 248402 218074 248582 218162
rect 248690 218074 248870 218162
rect 248978 218074 249158 218162
rect 249266 218074 249446 218162
rect 249554 218074 249734 218162
rect 249842 218074 250022 218162
rect 250130 218074 250310 218162
rect 250564 218074 250744 218162
rect 360436 218074 360560 218162
rect 360814 218074 360994 218162
rect 361102 218074 361282 218162
rect 361390 218074 361570 218162
rect 361678 218074 361858 218162
rect 361966 218074 362146 218162
rect 362254 218074 362434 218162
rect 362542 218074 362722 218162
rect 362830 218074 363010 218162
rect 363264 218074 363444 218162
rect 363552 218074 363732 218162
rect 363840 218074 364020 218162
rect 364128 218074 364308 218162
rect 364416 218074 364596 218162
rect 364704 218074 364884 218162
rect 364992 218074 365172 218162
rect 365280 218074 365460 218162
rect 365714 218074 365894 218162
rect 366002 218074 366182 218162
rect 366290 218074 366470 218162
rect 366578 218074 366758 218162
rect 366866 218074 367046 218162
rect 367154 218074 367334 218162
rect 367442 218074 367622 218162
rect 367730 218074 367910 218162
rect 243214 217598 243394 217686
rect 243502 217598 243682 217686
rect 243790 217598 243970 217686
rect 244078 217598 244258 217686
rect 244366 217598 244546 217686
rect 244654 217598 244834 217686
rect 244942 217598 245122 217686
rect 245230 217598 245410 217686
rect 245664 217598 245844 217686
rect 245952 217598 246132 217686
rect 246240 217598 246420 217686
rect 246528 217598 246708 217686
rect 246816 217598 246996 217686
rect 247104 217598 247284 217686
rect 247392 217598 247572 217686
rect 247680 217598 247860 217686
rect 248114 217598 248294 217686
rect 248402 217598 248582 217686
rect 248690 217598 248870 217686
rect 248978 217598 249158 217686
rect 249266 217598 249446 217686
rect 249554 217598 249734 217686
rect 249842 217598 250022 217686
rect 250130 217598 250310 217686
rect 250564 217598 250744 217686
rect 360436 217598 360560 217686
rect 360814 217598 360994 217686
rect 361102 217598 361282 217686
rect 361390 217598 361570 217686
rect 361678 217598 361858 217686
rect 361966 217598 362146 217686
rect 362254 217598 362434 217686
rect 362542 217598 362722 217686
rect 362830 217598 363010 217686
rect 363264 217598 363444 217686
rect 363552 217598 363732 217686
rect 363840 217598 364020 217686
rect 364128 217598 364308 217686
rect 364416 217598 364596 217686
rect 364704 217598 364884 217686
rect 364992 217598 365172 217686
rect 365280 217598 365460 217686
rect 365714 217598 365894 217686
rect 366002 217598 366182 217686
rect 366290 217598 366470 217686
rect 366578 217598 366758 217686
rect 366866 217598 367046 217686
rect 367154 217598 367334 217686
rect 367442 217598 367622 217686
rect 367730 217598 367910 217686
rect 243214 217382 243394 217470
rect 243502 217382 243682 217470
rect 243790 217382 243970 217470
rect 244078 217382 244258 217470
rect 244366 217382 244546 217470
rect 244654 217382 244834 217470
rect 244942 217382 245122 217470
rect 245230 217382 245410 217470
rect 245664 217382 245844 217470
rect 245952 217382 246132 217470
rect 246240 217382 246420 217470
rect 246528 217382 246708 217470
rect 246816 217382 246996 217470
rect 247104 217382 247284 217470
rect 247392 217382 247572 217470
rect 247680 217382 247860 217470
rect 248114 217382 248294 217470
rect 248402 217382 248582 217470
rect 248690 217382 248870 217470
rect 248978 217382 249158 217470
rect 249266 217382 249446 217470
rect 249554 217382 249734 217470
rect 249842 217382 250022 217470
rect 250130 217382 250310 217470
rect 250564 217382 250744 217470
rect 360436 217382 360560 217470
rect 360814 217382 360994 217470
rect 361102 217382 361282 217470
rect 361390 217382 361570 217470
rect 361678 217382 361858 217470
rect 361966 217382 362146 217470
rect 362254 217382 362434 217470
rect 362542 217382 362722 217470
rect 362830 217382 363010 217470
rect 363264 217382 363444 217470
rect 363552 217382 363732 217470
rect 363840 217382 364020 217470
rect 364128 217382 364308 217470
rect 364416 217382 364596 217470
rect 364704 217382 364884 217470
rect 364992 217382 365172 217470
rect 365280 217382 365460 217470
rect 365714 217382 365894 217470
rect 366002 217382 366182 217470
rect 366290 217382 366470 217470
rect 366578 217382 366758 217470
rect 366866 217382 367046 217470
rect 367154 217382 367334 217470
rect 367442 217382 367622 217470
rect 367730 217382 367910 217470
rect 243214 216906 243394 216994
rect 243502 216906 243682 216994
rect 243790 216906 243970 216994
rect 244078 216906 244258 216994
rect 244366 216906 244546 216994
rect 244654 216906 244834 216994
rect 244942 216906 245122 216994
rect 245230 216906 245410 216994
rect 245664 216906 245844 216994
rect 245952 216906 246132 216994
rect 246240 216906 246420 216994
rect 246528 216906 246708 216994
rect 246816 216906 246996 216994
rect 247104 216906 247284 216994
rect 247392 216906 247572 216994
rect 247680 216906 247860 216994
rect 248114 216906 248294 216994
rect 248402 216906 248582 216994
rect 248690 216906 248870 216994
rect 248978 216906 249158 216994
rect 249266 216906 249446 216994
rect 249554 216906 249734 216994
rect 249842 216906 250022 216994
rect 250130 216906 250310 216994
rect 250564 216906 250744 216994
rect 360436 216906 360560 216994
rect 360814 216906 360994 216994
rect 361102 216906 361282 216994
rect 361390 216906 361570 216994
rect 361678 216906 361858 216994
rect 361966 216906 362146 216994
rect 362254 216906 362434 216994
rect 362542 216906 362722 216994
rect 362830 216906 363010 216994
rect 363264 216906 363444 216994
rect 363552 216906 363732 216994
rect 363840 216906 364020 216994
rect 364128 216906 364308 216994
rect 364416 216906 364596 216994
rect 364704 216906 364884 216994
rect 364992 216906 365172 216994
rect 365280 216906 365460 216994
rect 365714 216906 365894 216994
rect 366002 216906 366182 216994
rect 366290 216906 366470 216994
rect 366578 216906 366758 216994
rect 366866 216906 367046 216994
rect 367154 216906 367334 216994
rect 367442 216906 367622 216994
rect 367730 216906 367910 216994
rect 243214 216690 243394 216778
rect 243502 216690 243682 216778
rect 243790 216690 243970 216778
rect 244078 216690 244258 216778
rect 244366 216690 244546 216778
rect 244654 216690 244834 216778
rect 244942 216690 245122 216778
rect 245230 216690 245410 216778
rect 245664 216690 245844 216778
rect 245952 216690 246132 216778
rect 246240 216690 246420 216778
rect 246528 216690 246708 216778
rect 246816 216690 246996 216778
rect 247104 216690 247284 216778
rect 247392 216690 247572 216778
rect 247680 216690 247860 216778
rect 248114 216690 248294 216778
rect 248402 216690 248582 216778
rect 248690 216690 248870 216778
rect 248978 216690 249158 216778
rect 249266 216690 249446 216778
rect 249554 216690 249734 216778
rect 249842 216690 250022 216778
rect 250130 216690 250310 216778
rect 250564 216690 250744 216778
rect 360436 216690 360560 216778
rect 360814 216690 360994 216778
rect 361102 216690 361282 216778
rect 361390 216690 361570 216778
rect 361678 216690 361858 216778
rect 361966 216690 362146 216778
rect 362254 216690 362434 216778
rect 362542 216690 362722 216778
rect 362830 216690 363010 216778
rect 363264 216690 363444 216778
rect 363552 216690 363732 216778
rect 363840 216690 364020 216778
rect 364128 216690 364308 216778
rect 364416 216690 364596 216778
rect 364704 216690 364884 216778
rect 364992 216690 365172 216778
rect 365280 216690 365460 216778
rect 365714 216690 365894 216778
rect 366002 216690 366182 216778
rect 366290 216690 366470 216778
rect 366578 216690 366758 216778
rect 366866 216690 367046 216778
rect 367154 216690 367334 216778
rect 367442 216690 367622 216778
rect 367730 216690 367910 216778
rect 243214 216214 243394 216302
rect 243502 216214 243682 216302
rect 243790 216214 243970 216302
rect 244078 216214 244258 216302
rect 244366 216214 244546 216302
rect 244654 216214 244834 216302
rect 244942 216214 245122 216302
rect 245230 216214 245410 216302
rect 245664 216214 245844 216302
rect 245952 216214 246132 216302
rect 246240 216214 246420 216302
rect 246528 216214 246708 216302
rect 246816 216214 246996 216302
rect 247104 216214 247284 216302
rect 247392 216214 247572 216302
rect 247680 216214 247860 216302
rect 248114 216214 248294 216302
rect 248402 216214 248582 216302
rect 248690 216214 248870 216302
rect 248978 216214 249158 216302
rect 249266 216214 249446 216302
rect 249554 216214 249734 216302
rect 249842 216214 250022 216302
rect 250130 216214 250310 216302
rect 250564 216214 250744 216302
rect 360436 216214 360560 216302
rect 360814 216214 360994 216302
rect 361102 216214 361282 216302
rect 361390 216214 361570 216302
rect 361678 216214 361858 216302
rect 361966 216214 362146 216302
rect 362254 216214 362434 216302
rect 362542 216214 362722 216302
rect 362830 216214 363010 216302
rect 363264 216214 363444 216302
rect 363552 216214 363732 216302
rect 363840 216214 364020 216302
rect 364128 216214 364308 216302
rect 364416 216214 364596 216302
rect 364704 216214 364884 216302
rect 364992 216214 365172 216302
rect 365280 216214 365460 216302
rect 365714 216214 365894 216302
rect 366002 216214 366182 216302
rect 366290 216214 366470 216302
rect 366578 216214 366758 216302
rect 366866 216214 367046 216302
rect 367154 216214 367334 216302
rect 367442 216214 367622 216302
rect 367730 216214 367910 216302
rect 243214 215998 243394 216086
rect 243502 215998 243682 216086
rect 243790 215998 243970 216086
rect 244078 215998 244258 216086
rect 244366 215998 244546 216086
rect 244654 215998 244834 216086
rect 244942 215998 245122 216086
rect 245230 215998 245410 216086
rect 245664 215998 245844 216086
rect 245952 215998 246132 216086
rect 246240 215998 246420 216086
rect 246528 215998 246708 216086
rect 246816 215998 246996 216086
rect 247104 215998 247284 216086
rect 247392 215998 247572 216086
rect 247680 215998 247860 216086
rect 248114 215998 248294 216086
rect 248402 215998 248582 216086
rect 248690 215998 248870 216086
rect 248978 215998 249158 216086
rect 249266 215998 249446 216086
rect 249554 215998 249734 216086
rect 249842 215998 250022 216086
rect 250130 215998 250310 216086
rect 250564 215998 250744 216086
rect 360436 215998 360560 216086
rect 360814 215998 360994 216086
rect 361102 215998 361282 216086
rect 361390 215998 361570 216086
rect 361678 215998 361858 216086
rect 361966 215998 362146 216086
rect 362254 215998 362434 216086
rect 362542 215998 362722 216086
rect 362830 215998 363010 216086
rect 363264 215998 363444 216086
rect 363552 215998 363732 216086
rect 363840 215998 364020 216086
rect 364128 215998 364308 216086
rect 364416 215998 364596 216086
rect 364704 215998 364884 216086
rect 364992 215998 365172 216086
rect 365280 215998 365460 216086
rect 365714 215998 365894 216086
rect 366002 215998 366182 216086
rect 366290 215998 366470 216086
rect 366578 215998 366758 216086
rect 366866 215998 367046 216086
rect 367154 215998 367334 216086
rect 367442 215998 367622 216086
rect 367730 215998 367910 216086
rect 243214 215522 243394 215610
rect 243502 215522 243682 215610
rect 243790 215522 243970 215610
rect 244078 215522 244258 215610
rect 244366 215522 244546 215610
rect 244654 215522 244834 215610
rect 244942 215522 245122 215610
rect 245230 215522 245410 215610
rect 245664 215522 245844 215610
rect 245952 215522 246132 215610
rect 246240 215522 246420 215610
rect 246528 215522 246708 215610
rect 246816 215522 246996 215610
rect 247104 215522 247284 215610
rect 247392 215522 247572 215610
rect 247680 215522 247860 215610
rect 248114 215522 248294 215610
rect 248402 215522 248582 215610
rect 248690 215522 248870 215610
rect 248978 215522 249158 215610
rect 249266 215522 249446 215610
rect 249554 215522 249734 215610
rect 249842 215522 250022 215610
rect 250130 215522 250310 215610
rect 250564 215522 250744 215610
rect 360436 215522 360560 215610
rect 360814 215522 360994 215610
rect 361102 215522 361282 215610
rect 361390 215522 361570 215610
rect 361678 215522 361858 215610
rect 361966 215522 362146 215610
rect 362254 215522 362434 215610
rect 362542 215522 362722 215610
rect 362830 215522 363010 215610
rect 363264 215522 363444 215610
rect 363552 215522 363732 215610
rect 363840 215522 364020 215610
rect 364128 215522 364308 215610
rect 364416 215522 364596 215610
rect 364704 215522 364884 215610
rect 364992 215522 365172 215610
rect 365280 215522 365460 215610
rect 365714 215522 365894 215610
rect 366002 215522 366182 215610
rect 366290 215522 366470 215610
rect 366578 215522 366758 215610
rect 366866 215522 367046 215610
rect 367154 215522 367334 215610
rect 367442 215522 367622 215610
rect 367730 215522 367910 215610
rect 243214 215048 243394 215136
rect 243502 215048 243682 215136
rect 243790 215048 243970 215136
rect 244078 215048 244258 215136
rect 244366 215048 244546 215136
rect 244654 215048 244834 215136
rect 244942 215048 245122 215136
rect 245230 215048 245410 215136
rect 245664 215048 245844 215136
rect 245952 215048 246132 215136
rect 246240 215048 246420 215136
rect 246528 215048 246708 215136
rect 246816 215048 246996 215136
rect 247104 215048 247284 215136
rect 247392 215048 247572 215136
rect 247680 215048 247860 215136
rect 248114 215048 248294 215136
rect 248402 215048 248582 215136
rect 248690 215048 248870 215136
rect 248978 215048 249158 215136
rect 249266 215048 249446 215136
rect 249554 215048 249734 215136
rect 249842 215048 250022 215136
rect 250130 215048 250310 215136
rect 250564 215048 250744 215136
rect 360436 215048 360560 215136
rect 360814 215048 360994 215136
rect 361102 215048 361282 215136
rect 361390 215048 361570 215136
rect 361678 215048 361858 215136
rect 361966 215048 362146 215136
rect 362254 215048 362434 215136
rect 362542 215048 362722 215136
rect 362830 215048 363010 215136
rect 363264 215048 363444 215136
rect 363552 215048 363732 215136
rect 363840 215048 364020 215136
rect 364128 215048 364308 215136
rect 364416 215048 364596 215136
rect 364704 215048 364884 215136
rect 364992 215048 365172 215136
rect 365280 215048 365460 215136
rect 365714 215048 365894 215136
rect 366002 215048 366182 215136
rect 366290 215048 366470 215136
rect 366578 215048 366758 215136
rect 366866 215048 367046 215136
rect 367154 215048 367334 215136
rect 367442 215048 367622 215136
rect 367730 215048 367910 215136
rect 243214 214572 243394 214660
rect 243502 214572 243682 214660
rect 243790 214572 243970 214660
rect 244078 214572 244258 214660
rect 244366 214572 244546 214660
rect 244654 214572 244834 214660
rect 244942 214572 245122 214660
rect 245230 214572 245410 214660
rect 245664 214572 245844 214660
rect 245952 214572 246132 214660
rect 246240 214572 246420 214660
rect 246528 214572 246708 214660
rect 246816 214572 246996 214660
rect 247104 214572 247284 214660
rect 247392 214572 247572 214660
rect 247680 214572 247860 214660
rect 248114 214572 248294 214660
rect 248402 214572 248582 214660
rect 248690 214572 248870 214660
rect 248978 214572 249158 214660
rect 249266 214572 249446 214660
rect 249554 214572 249734 214660
rect 249842 214572 250022 214660
rect 250130 214572 250310 214660
rect 250564 214572 250744 214660
rect 360436 214572 360560 214660
rect 360814 214572 360994 214660
rect 361102 214572 361282 214660
rect 361390 214572 361570 214660
rect 361678 214572 361858 214660
rect 361966 214572 362146 214660
rect 362254 214572 362434 214660
rect 362542 214572 362722 214660
rect 362830 214572 363010 214660
rect 363264 214572 363444 214660
rect 363552 214572 363732 214660
rect 363840 214572 364020 214660
rect 364128 214572 364308 214660
rect 364416 214572 364596 214660
rect 364704 214572 364884 214660
rect 364992 214572 365172 214660
rect 365280 214572 365460 214660
rect 365714 214572 365894 214660
rect 366002 214572 366182 214660
rect 366290 214572 366470 214660
rect 366578 214572 366758 214660
rect 366866 214572 367046 214660
rect 367154 214572 367334 214660
rect 367442 214572 367622 214660
rect 367730 214572 367910 214660
rect 243214 214356 243394 214444
rect 243502 214356 243682 214444
rect 243790 214356 243970 214444
rect 244078 214356 244258 214444
rect 244366 214356 244546 214444
rect 244654 214356 244834 214444
rect 244942 214356 245122 214444
rect 245230 214356 245410 214444
rect 245664 214356 245844 214444
rect 245952 214356 246132 214444
rect 246240 214356 246420 214444
rect 246528 214356 246708 214444
rect 246816 214356 246996 214444
rect 247104 214356 247284 214444
rect 247392 214356 247572 214444
rect 247680 214356 247860 214444
rect 248114 214356 248294 214444
rect 248402 214356 248582 214444
rect 248690 214356 248870 214444
rect 248978 214356 249158 214444
rect 249266 214356 249446 214444
rect 249554 214356 249734 214444
rect 249842 214356 250022 214444
rect 250130 214356 250310 214444
rect 250564 214356 250744 214444
rect 360436 214356 360560 214444
rect 360814 214356 360994 214444
rect 361102 214356 361282 214444
rect 361390 214356 361570 214444
rect 361678 214356 361858 214444
rect 361966 214356 362146 214444
rect 362254 214356 362434 214444
rect 362542 214356 362722 214444
rect 362830 214356 363010 214444
rect 363264 214356 363444 214444
rect 363552 214356 363732 214444
rect 363840 214356 364020 214444
rect 364128 214356 364308 214444
rect 364416 214356 364596 214444
rect 364704 214356 364884 214444
rect 364992 214356 365172 214444
rect 365280 214356 365460 214444
rect 365714 214356 365894 214444
rect 366002 214356 366182 214444
rect 366290 214356 366470 214444
rect 366578 214356 366758 214444
rect 366866 214356 367046 214444
rect 367154 214356 367334 214444
rect 367442 214356 367622 214444
rect 367730 214356 367910 214444
rect 243214 213880 243394 213968
rect 243502 213880 243682 213968
rect 243790 213880 243970 213968
rect 244078 213880 244258 213968
rect 244366 213880 244546 213968
rect 244654 213880 244834 213968
rect 244942 213880 245122 213968
rect 245230 213880 245410 213968
rect 245664 213880 245844 213968
rect 245952 213880 246132 213968
rect 246240 213880 246420 213968
rect 246528 213880 246708 213968
rect 246816 213880 246996 213968
rect 247104 213880 247284 213968
rect 247392 213880 247572 213968
rect 247680 213880 247860 213968
rect 248114 213880 248294 213968
rect 248402 213880 248582 213968
rect 248690 213880 248870 213968
rect 248978 213880 249158 213968
rect 249266 213880 249446 213968
rect 249554 213880 249734 213968
rect 249842 213880 250022 213968
rect 250130 213880 250310 213968
rect 250564 213880 250744 213968
rect 360436 213880 360560 213968
rect 360814 213880 360994 213968
rect 361102 213880 361282 213968
rect 361390 213880 361570 213968
rect 361678 213880 361858 213968
rect 361966 213880 362146 213968
rect 362254 213880 362434 213968
rect 362542 213880 362722 213968
rect 362830 213880 363010 213968
rect 363264 213880 363444 213968
rect 363552 213880 363732 213968
rect 363840 213880 364020 213968
rect 364128 213880 364308 213968
rect 364416 213880 364596 213968
rect 364704 213880 364884 213968
rect 364992 213880 365172 213968
rect 365280 213880 365460 213968
rect 365714 213880 365894 213968
rect 366002 213880 366182 213968
rect 366290 213880 366470 213968
rect 366578 213880 366758 213968
rect 366866 213880 367046 213968
rect 367154 213880 367334 213968
rect 367442 213880 367622 213968
rect 367730 213880 367910 213968
rect 243214 213664 243394 213752
rect 243502 213664 243682 213752
rect 243790 213664 243970 213752
rect 244078 213664 244258 213752
rect 244366 213664 244546 213752
rect 244654 213664 244834 213752
rect 244942 213664 245122 213752
rect 245230 213664 245410 213752
rect 245664 213664 245844 213752
rect 245952 213664 246132 213752
rect 246240 213664 246420 213752
rect 246528 213664 246708 213752
rect 246816 213664 246996 213752
rect 247104 213664 247284 213752
rect 247392 213664 247572 213752
rect 247680 213664 247860 213752
rect 248114 213664 248294 213752
rect 248402 213664 248582 213752
rect 248690 213664 248870 213752
rect 248978 213664 249158 213752
rect 249266 213664 249446 213752
rect 249554 213664 249734 213752
rect 249842 213664 250022 213752
rect 250130 213664 250310 213752
rect 250564 213664 250744 213752
rect 360436 213664 360560 213752
rect 360814 213664 360994 213752
rect 361102 213664 361282 213752
rect 361390 213664 361570 213752
rect 361678 213664 361858 213752
rect 361966 213664 362146 213752
rect 362254 213664 362434 213752
rect 362542 213664 362722 213752
rect 362830 213664 363010 213752
rect 363264 213664 363444 213752
rect 363552 213664 363732 213752
rect 363840 213664 364020 213752
rect 364128 213664 364308 213752
rect 364416 213664 364596 213752
rect 364704 213664 364884 213752
rect 364992 213664 365172 213752
rect 365280 213664 365460 213752
rect 365714 213664 365894 213752
rect 366002 213664 366182 213752
rect 366290 213664 366470 213752
rect 366578 213664 366758 213752
rect 366866 213664 367046 213752
rect 367154 213664 367334 213752
rect 367442 213664 367622 213752
rect 367730 213664 367910 213752
rect 243214 213188 243394 213276
rect 243502 213188 243682 213276
rect 243790 213188 243970 213276
rect 244078 213188 244258 213276
rect 244366 213188 244546 213276
rect 244654 213188 244834 213276
rect 244942 213188 245122 213276
rect 245230 213188 245410 213276
rect 245664 213188 245844 213276
rect 245952 213188 246132 213276
rect 246240 213188 246420 213276
rect 246528 213188 246708 213276
rect 246816 213188 246996 213276
rect 247104 213188 247284 213276
rect 247392 213188 247572 213276
rect 247680 213188 247860 213276
rect 248114 213188 248294 213276
rect 248402 213188 248582 213276
rect 248690 213188 248870 213276
rect 248978 213188 249158 213276
rect 249266 213188 249446 213276
rect 249554 213188 249734 213276
rect 249842 213188 250022 213276
rect 250130 213188 250310 213276
rect 250564 213188 250744 213276
rect 360436 213188 360560 213276
rect 360814 213188 360994 213276
rect 361102 213188 361282 213276
rect 361390 213188 361570 213276
rect 361678 213188 361858 213276
rect 361966 213188 362146 213276
rect 362254 213188 362434 213276
rect 362542 213188 362722 213276
rect 362830 213188 363010 213276
rect 363264 213188 363444 213276
rect 363552 213188 363732 213276
rect 363840 213188 364020 213276
rect 364128 213188 364308 213276
rect 364416 213188 364596 213276
rect 364704 213188 364884 213276
rect 364992 213188 365172 213276
rect 365280 213188 365460 213276
rect 365714 213188 365894 213276
rect 366002 213188 366182 213276
rect 366290 213188 366470 213276
rect 366578 213188 366758 213276
rect 366866 213188 367046 213276
rect 367154 213188 367334 213276
rect 367442 213188 367622 213276
rect 367730 213188 367910 213276
rect 243214 212972 243394 213060
rect 243502 212972 243682 213060
rect 243790 212972 243970 213060
rect 244078 212972 244258 213060
rect 244366 212972 244546 213060
rect 244654 212972 244834 213060
rect 244942 212972 245122 213060
rect 245230 212972 245410 213060
rect 245664 212972 245844 213060
rect 245952 212972 246132 213060
rect 246240 212972 246420 213060
rect 246528 212972 246708 213060
rect 246816 212972 246996 213060
rect 247104 212972 247284 213060
rect 247392 212972 247572 213060
rect 247680 212972 247860 213060
rect 248114 212972 248294 213060
rect 248402 212972 248582 213060
rect 248690 212972 248870 213060
rect 248978 212972 249158 213060
rect 249266 212972 249446 213060
rect 249554 212972 249734 213060
rect 249842 212972 250022 213060
rect 250130 212972 250310 213060
rect 250564 212972 250744 213060
rect 360436 212972 360560 213060
rect 360814 212972 360994 213060
rect 361102 212972 361282 213060
rect 361390 212972 361570 213060
rect 361678 212972 361858 213060
rect 361966 212972 362146 213060
rect 362254 212972 362434 213060
rect 362542 212972 362722 213060
rect 362830 212972 363010 213060
rect 363264 212972 363444 213060
rect 363552 212972 363732 213060
rect 363840 212972 364020 213060
rect 364128 212972 364308 213060
rect 364416 212972 364596 213060
rect 364704 212972 364884 213060
rect 364992 212972 365172 213060
rect 365280 212972 365460 213060
rect 365714 212972 365894 213060
rect 366002 212972 366182 213060
rect 366290 212972 366470 213060
rect 366578 212972 366758 213060
rect 366866 212972 367046 213060
rect 367154 212972 367334 213060
rect 367442 212972 367622 213060
rect 367730 212972 367910 213060
rect 243214 212496 243394 212584
rect 243502 212496 243682 212584
rect 243790 212496 243970 212584
rect 244078 212496 244258 212584
rect 244366 212496 244546 212584
rect 244654 212496 244834 212584
rect 244942 212496 245122 212584
rect 245230 212496 245410 212584
rect 245664 212496 245844 212584
rect 245952 212496 246132 212584
rect 246240 212496 246420 212584
rect 246528 212496 246708 212584
rect 246816 212496 246996 212584
rect 247104 212496 247284 212584
rect 247392 212496 247572 212584
rect 247680 212496 247860 212584
rect 248114 212496 248294 212584
rect 248402 212496 248582 212584
rect 248690 212496 248870 212584
rect 248978 212496 249158 212584
rect 249266 212496 249446 212584
rect 249554 212496 249734 212584
rect 249842 212496 250022 212584
rect 250130 212496 250310 212584
rect 250564 212496 250744 212584
rect 360436 212496 360560 212584
rect 360814 212496 360994 212584
rect 361102 212496 361282 212584
rect 361390 212496 361570 212584
rect 361678 212496 361858 212584
rect 361966 212496 362146 212584
rect 362254 212496 362434 212584
rect 362542 212496 362722 212584
rect 362830 212496 363010 212584
rect 363264 212496 363444 212584
rect 363552 212496 363732 212584
rect 363840 212496 364020 212584
rect 364128 212496 364308 212584
rect 364416 212496 364596 212584
rect 364704 212496 364884 212584
rect 364992 212496 365172 212584
rect 365280 212496 365460 212584
rect 365714 212496 365894 212584
rect 366002 212496 366182 212584
rect 366290 212496 366470 212584
rect 366578 212496 366758 212584
rect 366866 212496 367046 212584
rect 367154 212496 367334 212584
rect 367442 212496 367622 212584
rect 367730 212496 367910 212584
rect 243214 212022 243394 212110
rect 243502 212022 243682 212110
rect 243790 212022 243970 212110
rect 244078 212022 244258 212110
rect 244366 212022 244546 212110
rect 244654 212022 244834 212110
rect 244942 212022 245122 212110
rect 245230 212022 245410 212110
rect 245664 212022 245844 212110
rect 245952 212022 246132 212110
rect 246240 212022 246420 212110
rect 246528 212022 246708 212110
rect 246816 212022 246996 212110
rect 247104 212022 247284 212110
rect 247392 212022 247572 212110
rect 247680 212022 247860 212110
rect 248114 212022 248294 212110
rect 248402 212022 248582 212110
rect 248690 212022 248870 212110
rect 248978 212022 249158 212110
rect 249266 212022 249446 212110
rect 249554 212022 249734 212110
rect 249842 212022 250022 212110
rect 250130 212022 250310 212110
rect 250564 212022 250744 212110
rect 360436 212022 360560 212110
rect 360814 212022 360994 212110
rect 361102 212022 361282 212110
rect 361390 212022 361570 212110
rect 361678 212022 361858 212110
rect 361966 212022 362146 212110
rect 362254 212022 362434 212110
rect 362542 212022 362722 212110
rect 362830 212022 363010 212110
rect 363264 212022 363444 212110
rect 363552 212022 363732 212110
rect 363840 212022 364020 212110
rect 364128 212022 364308 212110
rect 364416 212022 364596 212110
rect 364704 212022 364884 212110
rect 364992 212022 365172 212110
rect 365280 212022 365460 212110
rect 365714 212022 365894 212110
rect 366002 212022 366182 212110
rect 366290 212022 366470 212110
rect 366578 212022 366758 212110
rect 366866 212022 367046 212110
rect 367154 212022 367334 212110
rect 367442 212022 367622 212110
rect 367730 212022 367910 212110
rect 243214 211546 243394 211634
rect 243502 211546 243682 211634
rect 243790 211546 243970 211634
rect 244078 211546 244258 211634
rect 244366 211546 244546 211634
rect 244654 211546 244834 211634
rect 244942 211546 245122 211634
rect 245230 211546 245410 211634
rect 245664 211546 245844 211634
rect 245952 211546 246132 211634
rect 246240 211546 246420 211634
rect 246528 211546 246708 211634
rect 246816 211546 246996 211634
rect 247104 211546 247284 211634
rect 247392 211546 247572 211634
rect 247680 211546 247860 211634
rect 248114 211546 248294 211634
rect 248402 211546 248582 211634
rect 248690 211546 248870 211634
rect 248978 211546 249158 211634
rect 249266 211546 249446 211634
rect 249554 211546 249734 211634
rect 249842 211546 250022 211634
rect 250130 211546 250310 211634
rect 250564 211546 250744 211634
rect 360436 211546 360560 211634
rect 360814 211546 360994 211634
rect 361102 211546 361282 211634
rect 361390 211546 361570 211634
rect 361678 211546 361858 211634
rect 361966 211546 362146 211634
rect 362254 211546 362434 211634
rect 362542 211546 362722 211634
rect 362830 211546 363010 211634
rect 363264 211546 363444 211634
rect 363552 211546 363732 211634
rect 363840 211546 364020 211634
rect 364128 211546 364308 211634
rect 364416 211546 364596 211634
rect 364704 211546 364884 211634
rect 364992 211546 365172 211634
rect 365280 211546 365460 211634
rect 365714 211546 365894 211634
rect 366002 211546 366182 211634
rect 366290 211546 366470 211634
rect 366578 211546 366758 211634
rect 366866 211546 367046 211634
rect 367154 211546 367334 211634
rect 367442 211546 367622 211634
rect 367730 211546 367910 211634
rect 243214 211330 243394 211418
rect 243502 211330 243682 211418
rect 243790 211330 243970 211418
rect 244078 211330 244258 211418
rect 244366 211330 244546 211418
rect 244654 211330 244834 211418
rect 244942 211330 245122 211418
rect 245230 211330 245410 211418
rect 245664 211330 245844 211418
rect 245952 211330 246132 211418
rect 246240 211330 246420 211418
rect 246528 211330 246708 211418
rect 246816 211330 246996 211418
rect 247104 211330 247284 211418
rect 247392 211330 247572 211418
rect 247680 211330 247860 211418
rect 248114 211330 248294 211418
rect 248402 211330 248582 211418
rect 248690 211330 248870 211418
rect 248978 211330 249158 211418
rect 249266 211330 249446 211418
rect 249554 211330 249734 211418
rect 249842 211330 250022 211418
rect 250130 211330 250310 211418
rect 250564 211330 250744 211418
rect 360436 211330 360560 211418
rect 360814 211330 360994 211418
rect 361102 211330 361282 211418
rect 361390 211330 361570 211418
rect 361678 211330 361858 211418
rect 361966 211330 362146 211418
rect 362254 211330 362434 211418
rect 362542 211330 362722 211418
rect 362830 211330 363010 211418
rect 363264 211330 363444 211418
rect 363552 211330 363732 211418
rect 363840 211330 364020 211418
rect 364128 211330 364308 211418
rect 364416 211330 364596 211418
rect 364704 211330 364884 211418
rect 364992 211330 365172 211418
rect 365280 211330 365460 211418
rect 365714 211330 365894 211418
rect 366002 211330 366182 211418
rect 366290 211330 366470 211418
rect 366578 211330 366758 211418
rect 366866 211330 367046 211418
rect 367154 211330 367334 211418
rect 367442 211330 367622 211418
rect 367730 211330 367910 211418
rect 243214 210854 243394 210942
rect 243502 210854 243682 210942
rect 243790 210854 243970 210942
rect 244078 210854 244258 210942
rect 244366 210854 244546 210942
rect 244654 210854 244834 210942
rect 244942 210854 245122 210942
rect 245230 210854 245410 210942
rect 245664 210854 245844 210942
rect 245952 210854 246132 210942
rect 246240 210854 246420 210942
rect 246528 210854 246708 210942
rect 246816 210854 246996 210942
rect 247104 210854 247284 210942
rect 247392 210854 247572 210942
rect 247680 210854 247860 210942
rect 248114 210854 248294 210942
rect 248402 210854 248582 210942
rect 248690 210854 248870 210942
rect 248978 210854 249158 210942
rect 249266 210854 249446 210942
rect 249554 210854 249734 210942
rect 249842 210854 250022 210942
rect 250130 210854 250310 210942
rect 250564 210854 250744 210942
rect 360436 210854 360560 210942
rect 360814 210854 360994 210942
rect 361102 210854 361282 210942
rect 361390 210854 361570 210942
rect 361678 210854 361858 210942
rect 361966 210854 362146 210942
rect 362254 210854 362434 210942
rect 362542 210854 362722 210942
rect 362830 210854 363010 210942
rect 363264 210854 363444 210942
rect 363552 210854 363732 210942
rect 363840 210854 364020 210942
rect 364128 210854 364308 210942
rect 364416 210854 364596 210942
rect 364704 210854 364884 210942
rect 364992 210854 365172 210942
rect 365280 210854 365460 210942
rect 365714 210854 365894 210942
rect 366002 210854 366182 210942
rect 366290 210854 366470 210942
rect 366578 210854 366758 210942
rect 366866 210854 367046 210942
rect 367154 210854 367334 210942
rect 367442 210854 367622 210942
rect 367730 210854 367910 210942
rect 243214 210638 243394 210726
rect 243502 210638 243682 210726
rect 243790 210638 243970 210726
rect 244078 210638 244258 210726
rect 244366 210638 244546 210726
rect 244654 210638 244834 210726
rect 244942 210638 245122 210726
rect 245230 210638 245410 210726
rect 245664 210638 245844 210726
rect 245952 210638 246132 210726
rect 246240 210638 246420 210726
rect 246528 210638 246708 210726
rect 246816 210638 246996 210726
rect 247104 210638 247284 210726
rect 247392 210638 247572 210726
rect 247680 210638 247860 210726
rect 248114 210638 248294 210726
rect 248402 210638 248582 210726
rect 248690 210638 248870 210726
rect 248978 210638 249158 210726
rect 249266 210638 249446 210726
rect 249554 210638 249734 210726
rect 249842 210638 250022 210726
rect 250130 210638 250310 210726
rect 250564 210638 250744 210726
rect 360436 210638 360560 210726
rect 360814 210638 360994 210726
rect 361102 210638 361282 210726
rect 361390 210638 361570 210726
rect 361678 210638 361858 210726
rect 361966 210638 362146 210726
rect 362254 210638 362434 210726
rect 362542 210638 362722 210726
rect 362830 210638 363010 210726
rect 363264 210638 363444 210726
rect 363552 210638 363732 210726
rect 363840 210638 364020 210726
rect 364128 210638 364308 210726
rect 364416 210638 364596 210726
rect 364704 210638 364884 210726
rect 364992 210638 365172 210726
rect 365280 210638 365460 210726
rect 365714 210638 365894 210726
rect 366002 210638 366182 210726
rect 366290 210638 366470 210726
rect 366578 210638 366758 210726
rect 366866 210638 367046 210726
rect 367154 210638 367334 210726
rect 367442 210638 367622 210726
rect 367730 210638 367910 210726
rect 243214 210162 243394 210250
rect 243502 210162 243682 210250
rect 243790 210162 243970 210250
rect 244078 210162 244258 210250
rect 244366 210162 244546 210250
rect 244654 210162 244834 210250
rect 244942 210162 245122 210250
rect 245230 210162 245410 210250
rect 245664 210162 245844 210250
rect 245952 210162 246132 210250
rect 246240 210162 246420 210250
rect 246528 210162 246708 210250
rect 246816 210162 246996 210250
rect 247104 210162 247284 210250
rect 247392 210162 247572 210250
rect 247680 210162 247860 210250
rect 248114 210162 248294 210250
rect 248402 210162 248582 210250
rect 248690 210162 248870 210250
rect 248978 210162 249158 210250
rect 249266 210162 249446 210250
rect 249554 210162 249734 210250
rect 249842 210162 250022 210250
rect 250130 210162 250310 210250
rect 250564 210162 250744 210250
rect 360436 210162 360560 210250
rect 360814 210162 360994 210250
rect 361102 210162 361282 210250
rect 361390 210162 361570 210250
rect 361678 210162 361858 210250
rect 361966 210162 362146 210250
rect 362254 210162 362434 210250
rect 362542 210162 362722 210250
rect 362830 210162 363010 210250
rect 363264 210162 363444 210250
rect 363552 210162 363732 210250
rect 363840 210162 364020 210250
rect 364128 210162 364308 210250
rect 364416 210162 364596 210250
rect 364704 210162 364884 210250
rect 364992 210162 365172 210250
rect 365280 210162 365460 210250
rect 365714 210162 365894 210250
rect 366002 210162 366182 210250
rect 366290 210162 366470 210250
rect 366578 210162 366758 210250
rect 366866 210162 367046 210250
rect 367154 210162 367334 210250
rect 367442 210162 367622 210250
rect 367730 210162 367910 210250
rect 243214 209946 243394 210034
rect 243502 209946 243682 210034
rect 243790 209946 243970 210034
rect 244078 209946 244258 210034
rect 244366 209946 244546 210034
rect 244654 209946 244834 210034
rect 244942 209946 245122 210034
rect 245230 209946 245410 210034
rect 245664 209946 245844 210034
rect 245952 209946 246132 210034
rect 246240 209946 246420 210034
rect 246528 209946 246708 210034
rect 246816 209946 246996 210034
rect 247104 209946 247284 210034
rect 247392 209946 247572 210034
rect 247680 209946 247860 210034
rect 248114 209946 248294 210034
rect 248402 209946 248582 210034
rect 248690 209946 248870 210034
rect 248978 209946 249158 210034
rect 249266 209946 249446 210034
rect 249554 209946 249734 210034
rect 249842 209946 250022 210034
rect 250130 209946 250310 210034
rect 250564 209946 250744 210034
rect 360436 209946 360560 210034
rect 360814 209946 360994 210034
rect 361102 209946 361282 210034
rect 361390 209946 361570 210034
rect 361678 209946 361858 210034
rect 361966 209946 362146 210034
rect 362254 209946 362434 210034
rect 362542 209946 362722 210034
rect 362830 209946 363010 210034
rect 363264 209946 363444 210034
rect 363552 209946 363732 210034
rect 363840 209946 364020 210034
rect 364128 209946 364308 210034
rect 364416 209946 364596 210034
rect 364704 209946 364884 210034
rect 364992 209946 365172 210034
rect 365280 209946 365460 210034
rect 365714 209946 365894 210034
rect 366002 209946 366182 210034
rect 366290 209946 366470 210034
rect 366578 209946 366758 210034
rect 366866 209946 367046 210034
rect 367154 209946 367334 210034
rect 367442 209946 367622 210034
rect 367730 209946 367910 210034
rect 243214 209470 243394 209558
rect 243502 209470 243682 209558
rect 243790 209470 243970 209558
rect 244078 209470 244258 209558
rect 244366 209470 244546 209558
rect 244654 209470 244834 209558
rect 244942 209470 245122 209558
rect 245230 209470 245410 209558
rect 245664 209470 245844 209558
rect 245952 209470 246132 209558
rect 246240 209470 246420 209558
rect 246528 209470 246708 209558
rect 246816 209470 246996 209558
rect 247104 209470 247284 209558
rect 247392 209470 247572 209558
rect 247680 209470 247860 209558
rect 248114 209470 248294 209558
rect 248402 209470 248582 209558
rect 248690 209470 248870 209558
rect 248978 209470 249158 209558
rect 249266 209470 249446 209558
rect 249554 209470 249734 209558
rect 249842 209470 250022 209558
rect 250130 209470 250310 209558
rect 250564 209470 250744 209558
rect 360436 209470 360560 209558
rect 360814 209470 360994 209558
rect 361102 209470 361282 209558
rect 361390 209470 361570 209558
rect 361678 209470 361858 209558
rect 361966 209470 362146 209558
rect 362254 209470 362434 209558
rect 362542 209470 362722 209558
rect 362830 209470 363010 209558
rect 363264 209470 363444 209558
rect 363552 209470 363732 209558
rect 363840 209470 364020 209558
rect 364128 209470 364308 209558
rect 364416 209470 364596 209558
rect 364704 209470 364884 209558
rect 364992 209470 365172 209558
rect 365280 209470 365460 209558
rect 365714 209470 365894 209558
rect 366002 209470 366182 209558
rect 366290 209470 366470 209558
rect 366578 209470 366758 209558
rect 366866 209470 367046 209558
rect 367154 209470 367334 209558
rect 367442 209470 367622 209558
rect 367730 209470 367910 209558
rect 243214 208996 243394 209084
rect 243502 208996 243682 209084
rect 243790 208996 243970 209084
rect 244078 208996 244258 209084
rect 244366 208996 244546 209084
rect 244654 208996 244834 209084
rect 244942 208996 245122 209084
rect 245230 208996 245410 209084
rect 245664 208996 245844 209084
rect 245952 208996 246132 209084
rect 246240 208996 246420 209084
rect 246528 208996 246708 209084
rect 246816 208996 246996 209084
rect 247104 208996 247284 209084
rect 247392 208996 247572 209084
rect 247680 208996 247860 209084
rect 248114 208996 248294 209084
rect 248402 208996 248582 209084
rect 248690 208996 248870 209084
rect 248978 208996 249158 209084
rect 249266 208996 249446 209084
rect 249554 208996 249734 209084
rect 249842 208996 250022 209084
rect 250130 208996 250310 209084
rect 250564 208996 250744 209084
rect 360436 208996 360560 209084
rect 360814 208996 360994 209084
rect 361102 208996 361282 209084
rect 361390 208996 361570 209084
rect 361678 208996 361858 209084
rect 361966 208996 362146 209084
rect 362254 208996 362434 209084
rect 362542 208996 362722 209084
rect 362830 208996 363010 209084
rect 363264 208996 363444 209084
rect 363552 208996 363732 209084
rect 363840 208996 364020 209084
rect 364128 208996 364308 209084
rect 364416 208996 364596 209084
rect 364704 208996 364884 209084
rect 364992 208996 365172 209084
rect 365280 208996 365460 209084
rect 365714 208996 365894 209084
rect 366002 208996 366182 209084
rect 366290 208996 366470 209084
rect 366578 208996 366758 209084
rect 366866 208996 367046 209084
rect 367154 208996 367334 209084
rect 367442 208996 367622 209084
rect 367730 208996 367910 209084
rect 243214 208520 243394 208608
rect 243502 208520 243682 208608
rect 243790 208520 243970 208608
rect 244078 208520 244258 208608
rect 244366 208520 244546 208608
rect 244654 208520 244834 208608
rect 244942 208520 245122 208608
rect 245230 208520 245410 208608
rect 245664 208520 245844 208608
rect 245952 208520 246132 208608
rect 246240 208520 246420 208608
rect 246528 208520 246708 208608
rect 246816 208520 246996 208608
rect 247104 208520 247284 208608
rect 247392 208520 247572 208608
rect 247680 208520 247860 208608
rect 248114 208520 248294 208608
rect 248402 208520 248582 208608
rect 248690 208520 248870 208608
rect 248978 208520 249158 208608
rect 249266 208520 249446 208608
rect 249554 208520 249734 208608
rect 249842 208520 250022 208608
rect 250130 208520 250310 208608
rect 250564 208520 250744 208608
rect 360436 208520 360560 208608
rect 360814 208520 360994 208608
rect 361102 208520 361282 208608
rect 361390 208520 361570 208608
rect 361678 208520 361858 208608
rect 361966 208520 362146 208608
rect 362254 208520 362434 208608
rect 362542 208520 362722 208608
rect 362830 208520 363010 208608
rect 363264 208520 363444 208608
rect 363552 208520 363732 208608
rect 363840 208520 364020 208608
rect 364128 208520 364308 208608
rect 364416 208520 364596 208608
rect 364704 208520 364884 208608
rect 364992 208520 365172 208608
rect 365280 208520 365460 208608
rect 365714 208520 365894 208608
rect 366002 208520 366182 208608
rect 366290 208520 366470 208608
rect 366578 208520 366758 208608
rect 366866 208520 367046 208608
rect 367154 208520 367334 208608
rect 367442 208520 367622 208608
rect 367730 208520 367910 208608
rect 243214 208304 243394 208392
rect 243502 208304 243682 208392
rect 243790 208304 243970 208392
rect 244078 208304 244258 208392
rect 244366 208304 244546 208392
rect 244654 208304 244834 208392
rect 244942 208304 245122 208392
rect 245230 208304 245410 208392
rect 245664 208304 245844 208392
rect 245952 208304 246132 208392
rect 246240 208304 246420 208392
rect 246528 208304 246708 208392
rect 246816 208304 246996 208392
rect 247104 208304 247284 208392
rect 247392 208304 247572 208392
rect 247680 208304 247860 208392
rect 248114 208304 248294 208392
rect 248402 208304 248582 208392
rect 248690 208304 248870 208392
rect 248978 208304 249158 208392
rect 249266 208304 249446 208392
rect 249554 208304 249734 208392
rect 249842 208304 250022 208392
rect 250130 208304 250310 208392
rect 250564 208304 250744 208392
rect 360436 208304 360560 208392
rect 360814 208304 360994 208392
rect 361102 208304 361282 208392
rect 361390 208304 361570 208392
rect 361678 208304 361858 208392
rect 361966 208304 362146 208392
rect 362254 208304 362434 208392
rect 362542 208304 362722 208392
rect 362830 208304 363010 208392
rect 363264 208304 363444 208392
rect 363552 208304 363732 208392
rect 363840 208304 364020 208392
rect 364128 208304 364308 208392
rect 364416 208304 364596 208392
rect 364704 208304 364884 208392
rect 364992 208304 365172 208392
rect 365280 208304 365460 208392
rect 365714 208304 365894 208392
rect 366002 208304 366182 208392
rect 366290 208304 366470 208392
rect 366578 208304 366758 208392
rect 366866 208304 367046 208392
rect 367154 208304 367334 208392
rect 367442 208304 367622 208392
rect 367730 208304 367910 208392
rect 243214 207828 243394 207916
rect 243502 207828 243682 207916
rect 243790 207828 243970 207916
rect 244078 207828 244258 207916
rect 244366 207828 244546 207916
rect 244654 207828 244834 207916
rect 244942 207828 245122 207916
rect 245230 207828 245410 207916
rect 245664 207828 245844 207916
rect 245952 207828 246132 207916
rect 246240 207828 246420 207916
rect 246528 207828 246708 207916
rect 246816 207828 246996 207916
rect 247104 207828 247284 207916
rect 247392 207828 247572 207916
rect 247680 207828 247860 207916
rect 248114 207828 248294 207916
rect 248402 207828 248582 207916
rect 248690 207828 248870 207916
rect 248978 207828 249158 207916
rect 249266 207828 249446 207916
rect 249554 207828 249734 207916
rect 249842 207828 250022 207916
rect 250130 207828 250310 207916
rect 250564 207828 250744 207916
rect 360436 207828 360560 207916
rect 360814 207828 360994 207916
rect 361102 207828 361282 207916
rect 361390 207828 361570 207916
rect 361678 207828 361858 207916
rect 361966 207828 362146 207916
rect 362254 207828 362434 207916
rect 362542 207828 362722 207916
rect 362830 207828 363010 207916
rect 363264 207828 363444 207916
rect 363552 207828 363732 207916
rect 363840 207828 364020 207916
rect 364128 207828 364308 207916
rect 364416 207828 364596 207916
rect 364704 207828 364884 207916
rect 364992 207828 365172 207916
rect 365280 207828 365460 207916
rect 365714 207828 365894 207916
rect 366002 207828 366182 207916
rect 366290 207828 366470 207916
rect 366578 207828 366758 207916
rect 366866 207828 367046 207916
rect 367154 207828 367334 207916
rect 367442 207828 367622 207916
rect 367730 207828 367910 207916
rect 243214 207612 243394 207700
rect 243502 207612 243682 207700
rect 243790 207612 243970 207700
rect 244078 207612 244258 207700
rect 244366 207612 244546 207700
rect 244654 207612 244834 207700
rect 244942 207612 245122 207700
rect 245230 207612 245410 207700
rect 245664 207612 245844 207700
rect 245952 207612 246132 207700
rect 246240 207612 246420 207700
rect 246528 207612 246708 207700
rect 246816 207612 246996 207700
rect 247104 207612 247284 207700
rect 247392 207612 247572 207700
rect 247680 207612 247860 207700
rect 248114 207612 248294 207700
rect 248402 207612 248582 207700
rect 248690 207612 248870 207700
rect 248978 207612 249158 207700
rect 249266 207612 249446 207700
rect 249554 207612 249734 207700
rect 249842 207612 250022 207700
rect 250130 207612 250310 207700
rect 250564 207612 250744 207700
rect 360436 207612 360560 207700
rect 360814 207612 360994 207700
rect 361102 207612 361282 207700
rect 361390 207612 361570 207700
rect 361678 207612 361858 207700
rect 361966 207612 362146 207700
rect 362254 207612 362434 207700
rect 362542 207612 362722 207700
rect 362830 207612 363010 207700
rect 363264 207612 363444 207700
rect 363552 207612 363732 207700
rect 363840 207612 364020 207700
rect 364128 207612 364308 207700
rect 364416 207612 364596 207700
rect 364704 207612 364884 207700
rect 364992 207612 365172 207700
rect 365280 207612 365460 207700
rect 365714 207612 365894 207700
rect 366002 207612 366182 207700
rect 366290 207612 366470 207700
rect 366578 207612 366758 207700
rect 366866 207612 367046 207700
rect 367154 207612 367334 207700
rect 367442 207612 367622 207700
rect 367730 207612 367910 207700
rect 243214 207136 243394 207224
rect 243502 207136 243682 207224
rect 243790 207136 243970 207224
rect 244078 207136 244258 207224
rect 244366 207136 244546 207224
rect 244654 207136 244834 207224
rect 244942 207136 245122 207224
rect 245230 207136 245410 207224
rect 245664 207136 245844 207224
rect 245952 207136 246132 207224
rect 246240 207136 246420 207224
rect 246528 207136 246708 207224
rect 246816 207136 246996 207224
rect 247104 207136 247284 207224
rect 247392 207136 247572 207224
rect 247680 207136 247860 207224
rect 248114 207136 248294 207224
rect 248402 207136 248582 207224
rect 248690 207136 248870 207224
rect 248978 207136 249158 207224
rect 249266 207136 249446 207224
rect 249554 207136 249734 207224
rect 249842 207136 250022 207224
rect 250130 207136 250310 207224
rect 250564 207136 250744 207224
rect 360436 207136 360560 207224
rect 360814 207136 360994 207224
rect 361102 207136 361282 207224
rect 361390 207136 361570 207224
rect 361678 207136 361858 207224
rect 361966 207136 362146 207224
rect 362254 207136 362434 207224
rect 362542 207136 362722 207224
rect 362830 207136 363010 207224
rect 363264 207136 363444 207224
rect 363552 207136 363732 207224
rect 363840 207136 364020 207224
rect 364128 207136 364308 207224
rect 364416 207136 364596 207224
rect 364704 207136 364884 207224
rect 364992 207136 365172 207224
rect 365280 207136 365460 207224
rect 365714 207136 365894 207224
rect 366002 207136 366182 207224
rect 366290 207136 366470 207224
rect 366578 207136 366758 207224
rect 366866 207136 367046 207224
rect 367154 207136 367334 207224
rect 367442 207136 367622 207224
rect 367730 207136 367910 207224
rect 243214 206920 243394 207008
rect 243502 206920 243682 207008
rect 243790 206920 243970 207008
rect 244078 206920 244258 207008
rect 244366 206920 244546 207008
rect 244654 206920 244834 207008
rect 244942 206920 245122 207008
rect 245230 206920 245410 207008
rect 245664 206920 245844 207008
rect 245952 206920 246132 207008
rect 246240 206920 246420 207008
rect 246528 206920 246708 207008
rect 246816 206920 246996 207008
rect 247104 206920 247284 207008
rect 247392 206920 247572 207008
rect 247680 206920 247860 207008
rect 248114 206920 248294 207008
rect 248402 206920 248582 207008
rect 248690 206920 248870 207008
rect 248978 206920 249158 207008
rect 249266 206920 249446 207008
rect 249554 206920 249734 207008
rect 249842 206920 250022 207008
rect 250130 206920 250310 207008
rect 250564 206920 250744 207008
rect 360436 206920 360560 207008
rect 360814 206920 360994 207008
rect 361102 206920 361282 207008
rect 361390 206920 361570 207008
rect 361678 206920 361858 207008
rect 361966 206920 362146 207008
rect 362254 206920 362434 207008
rect 362542 206920 362722 207008
rect 362830 206920 363010 207008
rect 363264 206920 363444 207008
rect 363552 206920 363732 207008
rect 363840 206920 364020 207008
rect 364128 206920 364308 207008
rect 364416 206920 364596 207008
rect 364704 206920 364884 207008
rect 364992 206920 365172 207008
rect 365280 206920 365460 207008
rect 365714 206920 365894 207008
rect 366002 206920 366182 207008
rect 366290 206920 366470 207008
rect 366578 206920 366758 207008
rect 366866 206920 367046 207008
rect 367154 206920 367334 207008
rect 367442 206920 367622 207008
rect 367730 206920 367910 207008
rect 243214 206444 243394 206532
rect 243502 206444 243682 206532
rect 243790 206444 243970 206532
rect 244078 206444 244258 206532
rect 244366 206444 244546 206532
rect 244654 206444 244834 206532
rect 244942 206444 245122 206532
rect 245230 206444 245410 206532
rect 245664 206444 245844 206532
rect 245952 206444 246132 206532
rect 246240 206444 246420 206532
rect 246528 206444 246708 206532
rect 246816 206444 246996 206532
rect 247104 206444 247284 206532
rect 247392 206444 247572 206532
rect 247680 206444 247860 206532
rect 248114 206444 248294 206532
rect 248402 206444 248582 206532
rect 248690 206444 248870 206532
rect 248978 206444 249158 206532
rect 249266 206444 249446 206532
rect 249554 206444 249734 206532
rect 249842 206444 250022 206532
rect 250130 206444 250310 206532
rect 250564 206444 250744 206532
rect 360436 206444 360560 206532
rect 360814 206444 360994 206532
rect 361102 206444 361282 206532
rect 361390 206444 361570 206532
rect 361678 206444 361858 206532
rect 361966 206444 362146 206532
rect 362254 206444 362434 206532
rect 362542 206444 362722 206532
rect 362830 206444 363010 206532
rect 363264 206444 363444 206532
rect 363552 206444 363732 206532
rect 363840 206444 364020 206532
rect 364128 206444 364308 206532
rect 364416 206444 364596 206532
rect 364704 206444 364884 206532
rect 364992 206444 365172 206532
rect 365280 206444 365460 206532
rect 365714 206444 365894 206532
rect 366002 206444 366182 206532
rect 366290 206444 366470 206532
rect 366578 206444 366758 206532
rect 366866 206444 367046 206532
rect 367154 206444 367334 206532
rect 367442 206444 367622 206532
rect 367730 206444 367910 206532
rect 243214 205970 243394 206058
rect 243502 205970 243682 206058
rect 243790 205970 243970 206058
rect 244078 205970 244258 206058
rect 244366 205970 244546 206058
rect 244654 205970 244834 206058
rect 244942 205970 245122 206058
rect 245230 205970 245410 206058
rect 245664 205970 245844 206058
rect 245952 205970 246132 206058
rect 246240 205970 246420 206058
rect 246528 205970 246708 206058
rect 246816 205970 246996 206058
rect 247104 205970 247284 206058
rect 247392 205970 247572 206058
rect 247680 205970 247860 206058
rect 248114 205970 248294 206058
rect 248402 205970 248582 206058
rect 248690 205970 248870 206058
rect 248978 205970 249158 206058
rect 249266 205970 249446 206058
rect 249554 205970 249734 206058
rect 249842 205970 250022 206058
rect 250130 205970 250310 206058
rect 250564 205970 250744 206058
rect 360436 205970 360560 206058
rect 360814 205970 360994 206058
rect 361102 205970 361282 206058
rect 361390 205970 361570 206058
rect 361678 205970 361858 206058
rect 361966 205970 362146 206058
rect 362254 205970 362434 206058
rect 362542 205970 362722 206058
rect 362830 205970 363010 206058
rect 363264 205970 363444 206058
rect 363552 205970 363732 206058
rect 363840 205970 364020 206058
rect 364128 205970 364308 206058
rect 364416 205970 364596 206058
rect 364704 205970 364884 206058
rect 364992 205970 365172 206058
rect 365280 205970 365460 206058
rect 365714 205970 365894 206058
rect 366002 205970 366182 206058
rect 366290 205970 366470 206058
rect 366578 205970 366758 206058
rect 366866 205970 367046 206058
rect 367154 205970 367334 206058
rect 367442 205970 367622 206058
rect 367730 205970 367910 206058
rect 243214 205494 243394 205582
rect 243502 205494 243682 205582
rect 243790 205494 243970 205582
rect 244078 205494 244258 205582
rect 244366 205494 244546 205582
rect 244654 205494 244834 205582
rect 244942 205494 245122 205582
rect 245230 205494 245410 205582
rect 245664 205494 245844 205582
rect 245952 205494 246132 205582
rect 246240 205494 246420 205582
rect 246528 205494 246708 205582
rect 246816 205494 246996 205582
rect 247104 205494 247284 205582
rect 247392 205494 247572 205582
rect 247680 205494 247860 205582
rect 248114 205494 248294 205582
rect 248402 205494 248582 205582
rect 248690 205494 248870 205582
rect 248978 205494 249158 205582
rect 249266 205494 249446 205582
rect 249554 205494 249734 205582
rect 249842 205494 250022 205582
rect 250130 205494 250310 205582
rect 250564 205494 250744 205582
rect 360436 205494 360560 205582
rect 360814 205494 360994 205582
rect 361102 205494 361282 205582
rect 361390 205494 361570 205582
rect 361678 205494 361858 205582
rect 361966 205494 362146 205582
rect 362254 205494 362434 205582
rect 362542 205494 362722 205582
rect 362830 205494 363010 205582
rect 363264 205494 363444 205582
rect 363552 205494 363732 205582
rect 363840 205494 364020 205582
rect 364128 205494 364308 205582
rect 364416 205494 364596 205582
rect 364704 205494 364884 205582
rect 364992 205494 365172 205582
rect 365280 205494 365460 205582
rect 365714 205494 365894 205582
rect 366002 205494 366182 205582
rect 366290 205494 366470 205582
rect 366578 205494 366758 205582
rect 366866 205494 367046 205582
rect 367154 205494 367334 205582
rect 367442 205494 367622 205582
rect 367730 205494 367910 205582
rect 243214 205278 243394 205366
rect 243502 205278 243682 205366
rect 243790 205278 243970 205366
rect 244078 205278 244258 205366
rect 244366 205278 244546 205366
rect 244654 205278 244834 205366
rect 244942 205278 245122 205366
rect 245230 205278 245410 205366
rect 245664 205278 245844 205366
rect 245952 205278 246132 205366
rect 246240 205278 246420 205366
rect 246528 205278 246708 205366
rect 246816 205278 246996 205366
rect 247104 205278 247284 205366
rect 247392 205278 247572 205366
rect 247680 205278 247860 205366
rect 248114 205278 248294 205366
rect 248402 205278 248582 205366
rect 248690 205278 248870 205366
rect 248978 205278 249158 205366
rect 249266 205278 249446 205366
rect 249554 205278 249734 205366
rect 249842 205278 250022 205366
rect 250130 205278 250310 205366
rect 250564 205278 250744 205366
rect 360436 205278 360560 205366
rect 360814 205278 360994 205366
rect 361102 205278 361282 205366
rect 361390 205278 361570 205366
rect 361678 205278 361858 205366
rect 361966 205278 362146 205366
rect 362254 205278 362434 205366
rect 362542 205278 362722 205366
rect 362830 205278 363010 205366
rect 363264 205278 363444 205366
rect 363552 205278 363732 205366
rect 363840 205278 364020 205366
rect 364128 205278 364308 205366
rect 364416 205278 364596 205366
rect 364704 205278 364884 205366
rect 364992 205278 365172 205366
rect 365280 205278 365460 205366
rect 365714 205278 365894 205366
rect 366002 205278 366182 205366
rect 366290 205278 366470 205366
rect 366578 205278 366758 205366
rect 366866 205278 367046 205366
rect 367154 205278 367334 205366
rect 367442 205278 367622 205366
rect 367730 205278 367910 205366
rect 243214 204802 243394 204890
rect 243502 204802 243682 204890
rect 243790 204802 243970 204890
rect 244078 204802 244258 204890
rect 244366 204802 244546 204890
rect 244654 204802 244834 204890
rect 244942 204802 245122 204890
rect 245230 204802 245410 204890
rect 245664 204802 245844 204890
rect 245952 204802 246132 204890
rect 246240 204802 246420 204890
rect 246528 204802 246708 204890
rect 246816 204802 246996 204890
rect 247104 204802 247284 204890
rect 247392 204802 247572 204890
rect 247680 204802 247860 204890
rect 248114 204802 248294 204890
rect 248402 204802 248582 204890
rect 248690 204802 248870 204890
rect 248978 204802 249158 204890
rect 249266 204802 249446 204890
rect 249554 204802 249734 204890
rect 249842 204802 250022 204890
rect 250130 204802 250310 204890
rect 250564 204802 250744 204890
rect 360436 204802 360560 204890
rect 360814 204802 360994 204890
rect 361102 204802 361282 204890
rect 361390 204802 361570 204890
rect 361678 204802 361858 204890
rect 361966 204802 362146 204890
rect 362254 204802 362434 204890
rect 362542 204802 362722 204890
rect 362830 204802 363010 204890
rect 363264 204802 363444 204890
rect 363552 204802 363732 204890
rect 363840 204802 364020 204890
rect 364128 204802 364308 204890
rect 364416 204802 364596 204890
rect 364704 204802 364884 204890
rect 364992 204802 365172 204890
rect 365280 204802 365460 204890
rect 365714 204802 365894 204890
rect 366002 204802 366182 204890
rect 366290 204802 366470 204890
rect 366578 204802 366758 204890
rect 366866 204802 367046 204890
rect 367154 204802 367334 204890
rect 367442 204802 367622 204890
rect 367730 204802 367910 204890
rect 243214 204586 243394 204674
rect 243502 204586 243682 204674
rect 243790 204586 243970 204674
rect 244078 204586 244258 204674
rect 244366 204586 244546 204674
rect 244654 204586 244834 204674
rect 244942 204586 245122 204674
rect 245230 204586 245410 204674
rect 245664 204586 245844 204674
rect 245952 204586 246132 204674
rect 246240 204586 246420 204674
rect 246528 204586 246708 204674
rect 246816 204586 246996 204674
rect 247104 204586 247284 204674
rect 247392 204586 247572 204674
rect 247680 204586 247860 204674
rect 248114 204586 248294 204674
rect 248402 204586 248582 204674
rect 248690 204586 248870 204674
rect 248978 204586 249158 204674
rect 249266 204586 249446 204674
rect 249554 204586 249734 204674
rect 249842 204586 250022 204674
rect 250130 204586 250310 204674
rect 250564 204586 250744 204674
rect 360436 204586 360560 204674
rect 360814 204586 360994 204674
rect 361102 204586 361282 204674
rect 361390 204586 361570 204674
rect 361678 204586 361858 204674
rect 361966 204586 362146 204674
rect 362254 204586 362434 204674
rect 362542 204586 362722 204674
rect 362830 204586 363010 204674
rect 363264 204586 363444 204674
rect 363552 204586 363732 204674
rect 363840 204586 364020 204674
rect 364128 204586 364308 204674
rect 364416 204586 364596 204674
rect 364704 204586 364884 204674
rect 364992 204586 365172 204674
rect 365280 204586 365460 204674
rect 365714 204586 365894 204674
rect 366002 204586 366182 204674
rect 366290 204586 366470 204674
rect 366578 204586 366758 204674
rect 366866 204586 367046 204674
rect 367154 204586 367334 204674
rect 367442 204586 367622 204674
rect 367730 204586 367910 204674
rect 243214 204110 243394 204198
rect 243502 204110 243682 204198
rect 243790 204110 243970 204198
rect 244078 204110 244258 204198
rect 244366 204110 244546 204198
rect 244654 204110 244834 204198
rect 244942 204110 245122 204198
rect 245230 204110 245410 204198
rect 245664 204110 245844 204198
rect 245952 204110 246132 204198
rect 246240 204110 246420 204198
rect 246528 204110 246708 204198
rect 246816 204110 246996 204198
rect 247104 204110 247284 204198
rect 247392 204110 247572 204198
rect 247680 204110 247860 204198
rect 248114 204110 248294 204198
rect 248402 204110 248582 204198
rect 248690 204110 248870 204198
rect 248978 204110 249158 204198
rect 249266 204110 249446 204198
rect 249554 204110 249734 204198
rect 249842 204110 250022 204198
rect 250130 204110 250310 204198
rect 250564 204110 250744 204198
rect 360436 204110 360560 204198
rect 360814 204110 360994 204198
rect 361102 204110 361282 204198
rect 361390 204110 361570 204198
rect 361678 204110 361858 204198
rect 361966 204110 362146 204198
rect 362254 204110 362434 204198
rect 362542 204110 362722 204198
rect 362830 204110 363010 204198
rect 363264 204110 363444 204198
rect 363552 204110 363732 204198
rect 363840 204110 364020 204198
rect 364128 204110 364308 204198
rect 364416 204110 364596 204198
rect 364704 204110 364884 204198
rect 364992 204110 365172 204198
rect 365280 204110 365460 204198
rect 365714 204110 365894 204198
rect 366002 204110 366182 204198
rect 366290 204110 366470 204198
rect 366578 204110 366758 204198
rect 366866 204110 367046 204198
rect 367154 204110 367334 204198
rect 367442 204110 367622 204198
rect 367730 204110 367910 204198
rect 243214 203894 243394 203982
rect 243502 203894 243682 203982
rect 243790 203894 243970 203982
rect 244078 203894 244258 203982
rect 244366 203894 244546 203982
rect 244654 203894 244834 203982
rect 244942 203894 245122 203982
rect 245230 203894 245410 203982
rect 245664 203894 245844 203982
rect 245952 203894 246132 203982
rect 246240 203894 246420 203982
rect 246528 203894 246708 203982
rect 246816 203894 246996 203982
rect 247104 203894 247284 203982
rect 247392 203894 247572 203982
rect 247680 203894 247860 203982
rect 248114 203894 248294 203982
rect 248402 203894 248582 203982
rect 248690 203894 248870 203982
rect 248978 203894 249158 203982
rect 249266 203894 249446 203982
rect 249554 203894 249734 203982
rect 249842 203894 250022 203982
rect 250130 203894 250310 203982
rect 250564 203894 250744 203982
rect 360436 203894 360560 203982
rect 360814 203894 360994 203982
rect 361102 203894 361282 203982
rect 361390 203894 361570 203982
rect 361678 203894 361858 203982
rect 361966 203894 362146 203982
rect 362254 203894 362434 203982
rect 362542 203894 362722 203982
rect 362830 203894 363010 203982
rect 363264 203894 363444 203982
rect 363552 203894 363732 203982
rect 363840 203894 364020 203982
rect 364128 203894 364308 203982
rect 364416 203894 364596 203982
rect 364704 203894 364884 203982
rect 364992 203894 365172 203982
rect 365280 203894 365460 203982
rect 365714 203894 365894 203982
rect 366002 203894 366182 203982
rect 366290 203894 366470 203982
rect 366578 203894 366758 203982
rect 366866 203894 367046 203982
rect 367154 203894 367334 203982
rect 367442 203894 367622 203982
rect 367730 203894 367910 203982
rect 243214 203418 243394 203506
rect 243502 203418 243682 203506
rect 243790 203418 243970 203506
rect 244078 203418 244258 203506
rect 244366 203418 244546 203506
rect 244654 203418 244834 203506
rect 244942 203418 245122 203506
rect 245230 203418 245410 203506
rect 245664 203418 245844 203506
rect 245952 203418 246132 203506
rect 246240 203418 246420 203506
rect 246528 203418 246708 203506
rect 246816 203418 246996 203506
rect 247104 203418 247284 203506
rect 247392 203418 247572 203506
rect 247680 203418 247860 203506
rect 248114 203418 248294 203506
rect 248402 203418 248582 203506
rect 248690 203418 248870 203506
rect 248978 203418 249158 203506
rect 249266 203418 249446 203506
rect 249554 203418 249734 203506
rect 249842 203418 250022 203506
rect 250130 203418 250310 203506
rect 250564 203418 250744 203506
rect 360436 203418 360560 203506
rect 360814 203418 360994 203506
rect 361102 203418 361282 203506
rect 361390 203418 361570 203506
rect 361678 203418 361858 203506
rect 361966 203418 362146 203506
rect 362254 203418 362434 203506
rect 362542 203418 362722 203506
rect 362830 203418 363010 203506
rect 363264 203418 363444 203506
rect 363552 203418 363732 203506
rect 363840 203418 364020 203506
rect 364128 203418 364308 203506
rect 364416 203418 364596 203506
rect 364704 203418 364884 203506
rect 364992 203418 365172 203506
rect 365280 203418 365460 203506
rect 365714 203418 365894 203506
rect 366002 203418 366182 203506
rect 366290 203418 366470 203506
rect 366578 203418 366758 203506
rect 366866 203418 367046 203506
rect 367154 203418 367334 203506
rect 367442 203418 367622 203506
rect 367730 203418 367910 203506
rect 243214 202944 243394 203032
rect 243502 202944 243682 203032
rect 243790 202944 243970 203032
rect 244078 202944 244258 203032
rect 244366 202944 244546 203032
rect 244654 202944 244834 203032
rect 244942 202944 245122 203032
rect 245230 202944 245410 203032
rect 245664 202944 245844 203032
rect 245952 202944 246132 203032
rect 246240 202944 246420 203032
rect 246528 202944 246708 203032
rect 246816 202944 246996 203032
rect 247104 202944 247284 203032
rect 247392 202944 247572 203032
rect 247680 202944 247860 203032
rect 248114 202944 248294 203032
rect 248402 202944 248582 203032
rect 248690 202944 248870 203032
rect 248978 202944 249158 203032
rect 249266 202944 249446 203032
rect 249554 202944 249734 203032
rect 249842 202944 250022 203032
rect 250130 202944 250310 203032
rect 250564 202944 250744 203032
rect 360436 202944 360560 203032
rect 360814 202944 360994 203032
rect 361102 202944 361282 203032
rect 361390 202944 361570 203032
rect 361678 202944 361858 203032
rect 361966 202944 362146 203032
rect 362254 202944 362434 203032
rect 362542 202944 362722 203032
rect 362830 202944 363010 203032
rect 363264 202944 363444 203032
rect 363552 202944 363732 203032
rect 363840 202944 364020 203032
rect 364128 202944 364308 203032
rect 364416 202944 364596 203032
rect 364704 202944 364884 203032
rect 364992 202944 365172 203032
rect 365280 202944 365460 203032
rect 365714 202944 365894 203032
rect 366002 202944 366182 203032
rect 366290 202944 366470 203032
rect 366578 202944 366758 203032
rect 366866 202944 367046 203032
rect 367154 202944 367334 203032
rect 367442 202944 367622 203032
rect 367730 202944 367910 203032
rect 243214 202468 243394 202556
rect 243502 202468 243682 202556
rect 243790 202468 243970 202556
rect 244078 202468 244258 202556
rect 244366 202468 244546 202556
rect 244654 202468 244834 202556
rect 244942 202468 245122 202556
rect 245230 202468 245410 202556
rect 245664 202468 245844 202556
rect 245952 202468 246132 202556
rect 246240 202468 246420 202556
rect 246528 202468 246708 202556
rect 246816 202468 246996 202556
rect 247104 202468 247284 202556
rect 247392 202468 247572 202556
rect 247680 202468 247860 202556
rect 248114 202468 248294 202556
rect 248402 202468 248582 202556
rect 248690 202468 248870 202556
rect 248978 202468 249158 202556
rect 249266 202468 249446 202556
rect 249554 202468 249734 202556
rect 249842 202468 250022 202556
rect 250130 202468 250310 202556
rect 250564 202468 250744 202556
rect 360436 202468 360560 202556
rect 360814 202468 360994 202556
rect 361102 202468 361282 202556
rect 361390 202468 361570 202556
rect 361678 202468 361858 202556
rect 361966 202468 362146 202556
rect 362254 202468 362434 202556
rect 362542 202468 362722 202556
rect 362830 202468 363010 202556
rect 363264 202468 363444 202556
rect 363552 202468 363732 202556
rect 363840 202468 364020 202556
rect 364128 202468 364308 202556
rect 364416 202468 364596 202556
rect 364704 202468 364884 202556
rect 364992 202468 365172 202556
rect 365280 202468 365460 202556
rect 365714 202468 365894 202556
rect 366002 202468 366182 202556
rect 366290 202468 366470 202556
rect 366578 202468 366758 202556
rect 366866 202468 367046 202556
rect 367154 202468 367334 202556
rect 367442 202468 367622 202556
rect 367730 202468 367910 202556
rect 243214 202252 243394 202340
rect 243502 202252 243682 202340
rect 243790 202252 243970 202340
rect 244078 202252 244258 202340
rect 244366 202252 244546 202340
rect 244654 202252 244834 202340
rect 244942 202252 245122 202340
rect 245230 202252 245410 202340
rect 245664 202252 245844 202340
rect 245952 202252 246132 202340
rect 246240 202252 246420 202340
rect 246528 202252 246708 202340
rect 246816 202252 246996 202340
rect 247104 202252 247284 202340
rect 247392 202252 247572 202340
rect 247680 202252 247860 202340
rect 248114 202252 248294 202340
rect 248402 202252 248582 202340
rect 248690 202252 248870 202340
rect 248978 202252 249158 202340
rect 249266 202252 249446 202340
rect 249554 202252 249734 202340
rect 249842 202252 250022 202340
rect 250130 202252 250310 202340
rect 250564 202252 250744 202340
rect 360436 202252 360560 202340
rect 360814 202252 360994 202340
rect 361102 202252 361282 202340
rect 361390 202252 361570 202340
rect 361678 202252 361858 202340
rect 361966 202252 362146 202340
rect 362254 202252 362434 202340
rect 362542 202252 362722 202340
rect 362830 202252 363010 202340
rect 363264 202252 363444 202340
rect 363552 202252 363732 202340
rect 363840 202252 364020 202340
rect 364128 202252 364308 202340
rect 364416 202252 364596 202340
rect 364704 202252 364884 202340
rect 364992 202252 365172 202340
rect 365280 202252 365460 202340
rect 365714 202252 365894 202340
rect 366002 202252 366182 202340
rect 366290 202252 366470 202340
rect 366578 202252 366758 202340
rect 366866 202252 367046 202340
rect 367154 202252 367334 202340
rect 367442 202252 367622 202340
rect 367730 202252 367910 202340
rect 243214 201776 243394 201864
rect 243502 201776 243682 201864
rect 243790 201776 243970 201864
rect 244078 201776 244258 201864
rect 244366 201776 244546 201864
rect 244654 201776 244834 201864
rect 244942 201776 245122 201864
rect 245230 201776 245410 201864
rect 245664 201776 245844 201864
rect 245952 201776 246132 201864
rect 246240 201776 246420 201864
rect 246528 201776 246708 201864
rect 246816 201776 246996 201864
rect 247104 201776 247284 201864
rect 247392 201776 247572 201864
rect 247680 201776 247860 201864
rect 248114 201776 248294 201864
rect 248402 201776 248582 201864
rect 248690 201776 248870 201864
rect 248978 201776 249158 201864
rect 249266 201776 249446 201864
rect 249554 201776 249734 201864
rect 249842 201776 250022 201864
rect 250130 201776 250310 201864
rect 250564 201776 250744 201864
rect 360436 201776 360560 201864
rect 360814 201776 360994 201864
rect 361102 201776 361282 201864
rect 361390 201776 361570 201864
rect 361678 201776 361858 201864
rect 361966 201776 362146 201864
rect 362254 201776 362434 201864
rect 362542 201776 362722 201864
rect 362830 201776 363010 201864
rect 363264 201776 363444 201864
rect 363552 201776 363732 201864
rect 363840 201776 364020 201864
rect 364128 201776 364308 201864
rect 364416 201776 364596 201864
rect 364704 201776 364884 201864
rect 364992 201776 365172 201864
rect 365280 201776 365460 201864
rect 365714 201776 365894 201864
rect 366002 201776 366182 201864
rect 366290 201776 366470 201864
rect 366578 201776 366758 201864
rect 366866 201776 367046 201864
rect 367154 201776 367334 201864
rect 367442 201776 367622 201864
rect 367730 201776 367910 201864
rect 243214 201560 243394 201648
rect 243502 201560 243682 201648
rect 243790 201560 243970 201648
rect 244078 201560 244258 201648
rect 244366 201560 244546 201648
rect 244654 201560 244834 201648
rect 244942 201560 245122 201648
rect 245230 201560 245410 201648
rect 245664 201560 245844 201648
rect 245952 201560 246132 201648
rect 246240 201560 246420 201648
rect 246528 201560 246708 201648
rect 246816 201560 246996 201648
rect 247104 201560 247284 201648
rect 247392 201560 247572 201648
rect 247680 201560 247860 201648
rect 248114 201560 248294 201648
rect 248402 201560 248582 201648
rect 248690 201560 248870 201648
rect 248978 201560 249158 201648
rect 249266 201560 249446 201648
rect 249554 201560 249734 201648
rect 249842 201560 250022 201648
rect 250130 201560 250310 201648
rect 250564 201560 250744 201648
rect 360436 201560 360560 201648
rect 360814 201560 360994 201648
rect 361102 201560 361282 201648
rect 361390 201560 361570 201648
rect 361678 201560 361858 201648
rect 361966 201560 362146 201648
rect 362254 201560 362434 201648
rect 362542 201560 362722 201648
rect 362830 201560 363010 201648
rect 363264 201560 363444 201648
rect 363552 201560 363732 201648
rect 363840 201560 364020 201648
rect 364128 201560 364308 201648
rect 364416 201560 364596 201648
rect 364704 201560 364884 201648
rect 364992 201560 365172 201648
rect 365280 201560 365460 201648
rect 365714 201560 365894 201648
rect 366002 201560 366182 201648
rect 366290 201560 366470 201648
rect 366578 201560 366758 201648
rect 366866 201560 367046 201648
rect 367154 201560 367334 201648
rect 367442 201560 367622 201648
rect 367730 201560 367910 201648
rect 243214 201084 243394 201172
rect 243502 201084 243682 201172
rect 243790 201084 243970 201172
rect 244078 201084 244258 201172
rect 244366 201084 244546 201172
rect 244654 201084 244834 201172
rect 244942 201084 245122 201172
rect 245230 201084 245410 201172
rect 245664 201084 245844 201172
rect 245952 201084 246132 201172
rect 246240 201084 246420 201172
rect 246528 201084 246708 201172
rect 246816 201084 246996 201172
rect 247104 201084 247284 201172
rect 247392 201084 247572 201172
rect 247680 201084 247860 201172
rect 248114 201084 248294 201172
rect 248402 201084 248582 201172
rect 248690 201084 248870 201172
rect 248978 201084 249158 201172
rect 249266 201084 249446 201172
rect 249554 201084 249734 201172
rect 249842 201084 250022 201172
rect 250130 201084 250310 201172
rect 250564 201084 250744 201172
rect 360436 201084 360560 201172
rect 360814 201084 360994 201172
rect 361102 201084 361282 201172
rect 361390 201084 361570 201172
rect 361678 201084 361858 201172
rect 361966 201084 362146 201172
rect 362254 201084 362434 201172
rect 362542 201084 362722 201172
rect 362830 201084 363010 201172
rect 363264 201084 363444 201172
rect 363552 201084 363732 201172
rect 363840 201084 364020 201172
rect 364128 201084 364308 201172
rect 364416 201084 364596 201172
rect 364704 201084 364884 201172
rect 364992 201084 365172 201172
rect 365280 201084 365460 201172
rect 365714 201084 365894 201172
rect 366002 201084 366182 201172
rect 366290 201084 366470 201172
rect 366578 201084 366758 201172
rect 366866 201084 367046 201172
rect 367154 201084 367334 201172
rect 367442 201084 367622 201172
rect 367730 201084 367910 201172
rect 243214 200868 243394 200956
rect 243502 200868 243682 200956
rect 243790 200868 243970 200956
rect 244078 200868 244258 200956
rect 244366 200868 244546 200956
rect 244654 200868 244834 200956
rect 244942 200868 245122 200956
rect 245230 200868 245410 200956
rect 245664 200868 245844 200956
rect 245952 200868 246132 200956
rect 246240 200868 246420 200956
rect 246528 200868 246708 200956
rect 246816 200868 246996 200956
rect 247104 200868 247284 200956
rect 247392 200868 247572 200956
rect 247680 200868 247860 200956
rect 248114 200868 248294 200956
rect 248402 200868 248582 200956
rect 248690 200868 248870 200956
rect 248978 200868 249158 200956
rect 249266 200868 249446 200956
rect 249554 200868 249734 200956
rect 249842 200868 250022 200956
rect 250130 200868 250310 200956
rect 250564 200868 250744 200956
rect 360436 200868 360560 200956
rect 360814 200868 360994 200956
rect 361102 200868 361282 200956
rect 361390 200868 361570 200956
rect 361678 200868 361858 200956
rect 361966 200868 362146 200956
rect 362254 200868 362434 200956
rect 362542 200868 362722 200956
rect 362830 200868 363010 200956
rect 363264 200868 363444 200956
rect 363552 200868 363732 200956
rect 363840 200868 364020 200956
rect 364128 200868 364308 200956
rect 364416 200868 364596 200956
rect 364704 200868 364884 200956
rect 364992 200868 365172 200956
rect 365280 200868 365460 200956
rect 365714 200868 365894 200956
rect 366002 200868 366182 200956
rect 366290 200868 366470 200956
rect 366578 200868 366758 200956
rect 366866 200868 367046 200956
rect 367154 200868 367334 200956
rect 367442 200868 367622 200956
rect 367730 200868 367910 200956
rect 243214 200392 243394 200480
rect 243502 200392 243682 200480
rect 243790 200392 243970 200480
rect 244078 200392 244258 200480
rect 244366 200392 244546 200480
rect 244654 200392 244834 200480
rect 244942 200392 245122 200480
rect 245230 200392 245410 200480
rect 245664 200392 245844 200480
rect 245952 200392 246132 200480
rect 246240 200392 246420 200480
rect 246528 200392 246708 200480
rect 246816 200392 246996 200480
rect 247104 200392 247284 200480
rect 247392 200392 247572 200480
rect 247680 200392 247860 200480
rect 248114 200392 248294 200480
rect 248402 200392 248582 200480
rect 248690 200392 248870 200480
rect 248978 200392 249158 200480
rect 249266 200392 249446 200480
rect 249554 200392 249734 200480
rect 249842 200392 250022 200480
rect 250130 200392 250310 200480
rect 250564 200392 250744 200480
rect 360436 200392 360560 200480
rect 360814 200392 360994 200480
rect 361102 200392 361282 200480
rect 361390 200392 361570 200480
rect 361678 200392 361858 200480
rect 361966 200392 362146 200480
rect 362254 200392 362434 200480
rect 362542 200392 362722 200480
rect 362830 200392 363010 200480
rect 363264 200392 363444 200480
rect 363552 200392 363732 200480
rect 363840 200392 364020 200480
rect 364128 200392 364308 200480
rect 364416 200392 364596 200480
rect 364704 200392 364884 200480
rect 364992 200392 365172 200480
rect 365280 200392 365460 200480
rect 365714 200392 365894 200480
rect 366002 200392 366182 200480
rect 366290 200392 366470 200480
rect 366578 200392 366758 200480
rect 366866 200392 367046 200480
rect 367154 200392 367334 200480
rect 367442 200392 367622 200480
rect 367730 200392 367910 200480
rect 243214 199918 243394 200006
rect 243502 199918 243682 200006
rect 243790 199918 243970 200006
rect 244078 199918 244258 200006
rect 244366 199918 244546 200006
rect 244654 199918 244834 200006
rect 244942 199918 245122 200006
rect 245230 199918 245410 200006
rect 245664 199918 245844 200006
rect 245952 199918 246132 200006
rect 246240 199918 246420 200006
rect 246528 199918 246708 200006
rect 246816 199918 246996 200006
rect 247104 199918 247284 200006
rect 247392 199918 247572 200006
rect 247680 199918 247860 200006
rect 248114 199918 248294 200006
rect 248402 199918 248582 200006
rect 248690 199918 248870 200006
rect 248978 199918 249158 200006
rect 249266 199918 249446 200006
rect 249554 199918 249734 200006
rect 249842 199918 250022 200006
rect 250130 199918 250310 200006
rect 250564 199918 250744 200006
rect 360436 199918 360560 200006
rect 360814 199918 360994 200006
rect 361102 199918 361282 200006
rect 361390 199918 361570 200006
rect 361678 199918 361858 200006
rect 361966 199918 362146 200006
rect 362254 199918 362434 200006
rect 362542 199918 362722 200006
rect 362830 199918 363010 200006
rect 363264 199918 363444 200006
rect 363552 199918 363732 200006
rect 363840 199918 364020 200006
rect 364128 199918 364308 200006
rect 364416 199918 364596 200006
rect 364704 199918 364884 200006
rect 364992 199918 365172 200006
rect 365280 199918 365460 200006
rect 365714 199918 365894 200006
rect 366002 199918 366182 200006
rect 366290 199918 366470 200006
rect 366578 199918 366758 200006
rect 366866 199918 367046 200006
rect 367154 199918 367334 200006
rect 367442 199918 367622 200006
rect 367730 199918 367910 200006
rect 243214 199442 243394 199530
rect 243502 199442 243682 199530
rect 243790 199442 243970 199530
rect 244078 199442 244258 199530
rect 244366 199442 244546 199530
rect 244654 199442 244834 199530
rect 244942 199442 245122 199530
rect 245230 199442 245410 199530
rect 245664 199442 245844 199530
rect 245952 199442 246132 199530
rect 246240 199442 246420 199530
rect 246528 199442 246708 199530
rect 246816 199442 246996 199530
rect 247104 199442 247284 199530
rect 247392 199442 247572 199530
rect 247680 199442 247860 199530
rect 248114 199442 248294 199530
rect 248402 199442 248582 199530
rect 248690 199442 248870 199530
rect 248978 199442 249158 199530
rect 249266 199442 249446 199530
rect 249554 199442 249734 199530
rect 249842 199442 250022 199530
rect 250130 199442 250310 199530
rect 250564 199442 250744 199530
rect 360436 199442 360560 199530
rect 360814 199442 360994 199530
rect 361102 199442 361282 199530
rect 361390 199442 361570 199530
rect 361678 199442 361858 199530
rect 361966 199442 362146 199530
rect 362254 199442 362434 199530
rect 362542 199442 362722 199530
rect 362830 199442 363010 199530
rect 363264 199442 363444 199530
rect 363552 199442 363732 199530
rect 363840 199442 364020 199530
rect 364128 199442 364308 199530
rect 364416 199442 364596 199530
rect 364704 199442 364884 199530
rect 364992 199442 365172 199530
rect 365280 199442 365460 199530
rect 365714 199442 365894 199530
rect 366002 199442 366182 199530
rect 366290 199442 366470 199530
rect 366578 199442 366758 199530
rect 366866 199442 367046 199530
rect 367154 199442 367334 199530
rect 367442 199442 367622 199530
rect 367730 199442 367910 199530
rect 243214 199226 243394 199314
rect 243502 199226 243682 199314
rect 243790 199226 243970 199314
rect 244078 199226 244258 199314
rect 244366 199226 244546 199314
rect 244654 199226 244834 199314
rect 244942 199226 245122 199314
rect 245230 199226 245410 199314
rect 245664 199226 245844 199314
rect 245952 199226 246132 199314
rect 246240 199226 246420 199314
rect 246528 199226 246708 199314
rect 246816 199226 246996 199314
rect 247104 199226 247284 199314
rect 247392 199226 247572 199314
rect 247680 199226 247860 199314
rect 248114 199226 248294 199314
rect 248402 199226 248582 199314
rect 248690 199226 248870 199314
rect 248978 199226 249158 199314
rect 249266 199226 249446 199314
rect 249554 199226 249734 199314
rect 249842 199226 250022 199314
rect 250130 199226 250310 199314
rect 250564 199226 250744 199314
rect 360436 199226 360560 199314
rect 360814 199226 360994 199314
rect 361102 199226 361282 199314
rect 361390 199226 361570 199314
rect 361678 199226 361858 199314
rect 361966 199226 362146 199314
rect 362254 199226 362434 199314
rect 362542 199226 362722 199314
rect 362830 199226 363010 199314
rect 363264 199226 363444 199314
rect 363552 199226 363732 199314
rect 363840 199226 364020 199314
rect 364128 199226 364308 199314
rect 364416 199226 364596 199314
rect 364704 199226 364884 199314
rect 364992 199226 365172 199314
rect 365280 199226 365460 199314
rect 365714 199226 365894 199314
rect 366002 199226 366182 199314
rect 366290 199226 366470 199314
rect 366578 199226 366758 199314
rect 366866 199226 367046 199314
rect 367154 199226 367334 199314
rect 367442 199226 367622 199314
rect 367730 199226 367910 199314
rect 243214 198750 243394 198838
rect 243502 198750 243682 198838
rect 243790 198750 243970 198838
rect 244078 198750 244258 198838
rect 244366 198750 244546 198838
rect 244654 198750 244834 198838
rect 244942 198750 245122 198838
rect 245230 198750 245410 198838
rect 245664 198750 245844 198838
rect 245952 198750 246132 198838
rect 246240 198750 246420 198838
rect 246528 198750 246708 198838
rect 246816 198750 246996 198838
rect 247104 198750 247284 198838
rect 247392 198750 247572 198838
rect 247680 198750 247860 198838
rect 248114 198750 248294 198838
rect 248402 198750 248582 198838
rect 248690 198750 248870 198838
rect 248978 198750 249158 198838
rect 249266 198750 249446 198838
rect 249554 198750 249734 198838
rect 249842 198750 250022 198838
rect 250130 198750 250310 198838
rect 250564 198750 250744 198838
rect 360436 198750 360560 198838
rect 360814 198750 360994 198838
rect 361102 198750 361282 198838
rect 361390 198750 361570 198838
rect 361678 198750 361858 198838
rect 361966 198750 362146 198838
rect 362254 198750 362434 198838
rect 362542 198750 362722 198838
rect 362830 198750 363010 198838
rect 363264 198750 363444 198838
rect 363552 198750 363732 198838
rect 363840 198750 364020 198838
rect 364128 198750 364308 198838
rect 364416 198750 364596 198838
rect 364704 198750 364884 198838
rect 364992 198750 365172 198838
rect 365280 198750 365460 198838
rect 365714 198750 365894 198838
rect 366002 198750 366182 198838
rect 366290 198750 366470 198838
rect 366578 198750 366758 198838
rect 366866 198750 367046 198838
rect 367154 198750 367334 198838
rect 367442 198750 367622 198838
rect 367730 198750 367910 198838
rect 243214 198534 243394 198622
rect 243502 198534 243682 198622
rect 243790 198534 243970 198622
rect 244078 198534 244258 198622
rect 244366 198534 244546 198622
rect 244654 198534 244834 198622
rect 244942 198534 245122 198622
rect 245230 198534 245410 198622
rect 245664 198534 245844 198622
rect 245952 198534 246132 198622
rect 246240 198534 246420 198622
rect 246528 198534 246708 198622
rect 246816 198534 246996 198622
rect 247104 198534 247284 198622
rect 247392 198534 247572 198622
rect 247680 198534 247860 198622
rect 248114 198534 248294 198622
rect 248402 198534 248582 198622
rect 248690 198534 248870 198622
rect 248978 198534 249158 198622
rect 249266 198534 249446 198622
rect 249554 198534 249734 198622
rect 249842 198534 250022 198622
rect 250130 198534 250310 198622
rect 250564 198534 250744 198622
rect 360436 198534 360560 198622
rect 360814 198534 360994 198622
rect 361102 198534 361282 198622
rect 361390 198534 361570 198622
rect 361678 198534 361858 198622
rect 361966 198534 362146 198622
rect 362254 198534 362434 198622
rect 362542 198534 362722 198622
rect 362830 198534 363010 198622
rect 363264 198534 363444 198622
rect 363552 198534 363732 198622
rect 363840 198534 364020 198622
rect 364128 198534 364308 198622
rect 364416 198534 364596 198622
rect 364704 198534 364884 198622
rect 364992 198534 365172 198622
rect 365280 198534 365460 198622
rect 365714 198534 365894 198622
rect 366002 198534 366182 198622
rect 366290 198534 366470 198622
rect 366578 198534 366758 198622
rect 366866 198534 367046 198622
rect 367154 198534 367334 198622
rect 367442 198534 367622 198622
rect 367730 198534 367910 198622
rect 243214 198058 243394 198146
rect 243502 198058 243682 198146
rect 243790 198058 243970 198146
rect 244078 198058 244258 198146
rect 244366 198058 244546 198146
rect 244654 198058 244834 198146
rect 244942 198058 245122 198146
rect 245230 198058 245410 198146
rect 245664 198058 245844 198146
rect 245952 198058 246132 198146
rect 246240 198058 246420 198146
rect 246528 198058 246708 198146
rect 246816 198058 246996 198146
rect 247104 198058 247284 198146
rect 247392 198058 247572 198146
rect 247680 198058 247860 198146
rect 248114 198058 248294 198146
rect 248402 198058 248582 198146
rect 248690 198058 248870 198146
rect 248978 198058 249158 198146
rect 249266 198058 249446 198146
rect 249554 198058 249734 198146
rect 249842 198058 250022 198146
rect 250130 198058 250310 198146
rect 250564 198058 250744 198146
rect 360436 198058 360560 198146
rect 360814 198058 360994 198146
rect 361102 198058 361282 198146
rect 361390 198058 361570 198146
rect 361678 198058 361858 198146
rect 361966 198058 362146 198146
rect 362254 198058 362434 198146
rect 362542 198058 362722 198146
rect 362830 198058 363010 198146
rect 363264 198058 363444 198146
rect 363552 198058 363732 198146
rect 363840 198058 364020 198146
rect 364128 198058 364308 198146
rect 364416 198058 364596 198146
rect 364704 198058 364884 198146
rect 364992 198058 365172 198146
rect 365280 198058 365460 198146
rect 365714 198058 365894 198146
rect 366002 198058 366182 198146
rect 366290 198058 366470 198146
rect 366578 198058 366758 198146
rect 366866 198058 367046 198146
rect 367154 198058 367334 198146
rect 367442 198058 367622 198146
rect 367730 198058 367910 198146
rect 243214 197842 243394 197930
rect 243502 197842 243682 197930
rect 243790 197842 243970 197930
rect 244078 197842 244258 197930
rect 244366 197842 244546 197930
rect 244654 197842 244834 197930
rect 244942 197842 245122 197930
rect 245230 197842 245410 197930
rect 245664 197842 245844 197930
rect 245952 197842 246132 197930
rect 246240 197842 246420 197930
rect 246528 197842 246708 197930
rect 246816 197842 246996 197930
rect 247104 197842 247284 197930
rect 247392 197842 247572 197930
rect 247680 197842 247860 197930
rect 248114 197842 248294 197930
rect 248402 197842 248582 197930
rect 248690 197842 248870 197930
rect 248978 197842 249158 197930
rect 249266 197842 249446 197930
rect 249554 197842 249734 197930
rect 249842 197842 250022 197930
rect 250130 197842 250310 197930
rect 250564 197842 250744 197930
rect 360436 197842 360560 197930
rect 360814 197842 360994 197930
rect 361102 197842 361282 197930
rect 361390 197842 361570 197930
rect 361678 197842 361858 197930
rect 361966 197842 362146 197930
rect 362254 197842 362434 197930
rect 362542 197842 362722 197930
rect 362830 197842 363010 197930
rect 363264 197842 363444 197930
rect 363552 197842 363732 197930
rect 363840 197842 364020 197930
rect 364128 197842 364308 197930
rect 364416 197842 364596 197930
rect 364704 197842 364884 197930
rect 364992 197842 365172 197930
rect 365280 197842 365460 197930
rect 365714 197842 365894 197930
rect 366002 197842 366182 197930
rect 366290 197842 366470 197930
rect 366578 197842 366758 197930
rect 366866 197842 367046 197930
rect 367154 197842 367334 197930
rect 367442 197842 367622 197930
rect 367730 197842 367910 197930
rect 243214 197366 243394 197454
rect 243502 197366 243682 197454
rect 243790 197366 243970 197454
rect 244078 197366 244258 197454
rect 244366 197366 244546 197454
rect 244654 197366 244834 197454
rect 244942 197366 245122 197454
rect 245230 197366 245410 197454
rect 245664 197366 245844 197454
rect 245952 197366 246132 197454
rect 246240 197366 246420 197454
rect 246528 197366 246708 197454
rect 246816 197366 246996 197454
rect 247104 197366 247284 197454
rect 247392 197366 247572 197454
rect 247680 197366 247860 197454
rect 248114 197366 248294 197454
rect 248402 197366 248582 197454
rect 248690 197366 248870 197454
rect 248978 197366 249158 197454
rect 249266 197366 249446 197454
rect 249554 197366 249734 197454
rect 249842 197366 250022 197454
rect 250130 197366 250310 197454
rect 250564 197366 250744 197454
rect 360436 197366 360560 197454
rect 360814 197366 360994 197454
rect 361102 197366 361282 197454
rect 361390 197366 361570 197454
rect 361678 197366 361858 197454
rect 361966 197366 362146 197454
rect 362254 197366 362434 197454
rect 362542 197366 362722 197454
rect 362830 197366 363010 197454
rect 363264 197366 363444 197454
rect 363552 197366 363732 197454
rect 363840 197366 364020 197454
rect 364128 197366 364308 197454
rect 364416 197366 364596 197454
rect 364704 197366 364884 197454
rect 364992 197366 365172 197454
rect 365280 197366 365460 197454
rect 365714 197366 365894 197454
rect 366002 197366 366182 197454
rect 366290 197366 366470 197454
rect 366578 197366 366758 197454
rect 366866 197366 367046 197454
rect 367154 197366 367334 197454
rect 367442 197366 367622 197454
rect 367730 197366 367910 197454
rect 243214 196892 243394 196980
rect 243502 196892 243682 196980
rect 243790 196892 243970 196980
rect 244078 196892 244258 196980
rect 244366 196892 244546 196980
rect 244654 196892 244834 196980
rect 244942 196892 245122 196980
rect 245230 196892 245410 196980
rect 245664 196892 245844 196980
rect 245952 196892 246132 196980
rect 246240 196892 246420 196980
rect 246528 196892 246708 196980
rect 246816 196892 246996 196980
rect 247104 196892 247284 196980
rect 247392 196892 247572 196980
rect 247680 196892 247860 196980
rect 248114 196892 248294 196980
rect 248402 196892 248582 196980
rect 248690 196892 248870 196980
rect 248978 196892 249158 196980
rect 249266 196892 249446 196980
rect 249554 196892 249734 196980
rect 249842 196892 250022 196980
rect 250130 196892 250310 196980
rect 250564 196892 250744 196980
rect 360436 196892 360560 196980
rect 360814 196892 360994 196980
rect 361102 196892 361282 196980
rect 361390 196892 361570 196980
rect 361678 196892 361858 196980
rect 361966 196892 362146 196980
rect 362254 196892 362434 196980
rect 362542 196892 362722 196980
rect 362830 196892 363010 196980
rect 363264 196892 363444 196980
rect 363552 196892 363732 196980
rect 363840 196892 364020 196980
rect 364128 196892 364308 196980
rect 364416 196892 364596 196980
rect 364704 196892 364884 196980
rect 364992 196892 365172 196980
rect 365280 196892 365460 196980
rect 365714 196892 365894 196980
rect 366002 196892 366182 196980
rect 366290 196892 366470 196980
rect 366578 196892 366758 196980
rect 366866 196892 367046 196980
rect 367154 196892 367334 196980
rect 367442 196892 367622 196980
rect 367730 196892 367910 196980
rect 243214 196416 243394 196504
rect 243502 196416 243682 196504
rect 243790 196416 243970 196504
rect 244078 196416 244258 196504
rect 244366 196416 244546 196504
rect 244654 196416 244834 196504
rect 244942 196416 245122 196504
rect 245230 196416 245410 196504
rect 245664 196416 245844 196504
rect 245952 196416 246132 196504
rect 246240 196416 246420 196504
rect 246528 196416 246708 196504
rect 246816 196416 246996 196504
rect 247104 196416 247284 196504
rect 247392 196416 247572 196504
rect 247680 196416 247860 196504
rect 248114 196416 248294 196504
rect 248402 196416 248582 196504
rect 248690 196416 248870 196504
rect 248978 196416 249158 196504
rect 249266 196416 249446 196504
rect 249554 196416 249734 196504
rect 249842 196416 250022 196504
rect 250130 196416 250310 196504
rect 250564 196416 250744 196504
rect 360436 196416 360560 196504
rect 360814 196416 360994 196504
rect 361102 196416 361282 196504
rect 361390 196416 361570 196504
rect 361678 196416 361858 196504
rect 361966 196416 362146 196504
rect 362254 196416 362434 196504
rect 362542 196416 362722 196504
rect 362830 196416 363010 196504
rect 363264 196416 363444 196504
rect 363552 196416 363732 196504
rect 363840 196416 364020 196504
rect 364128 196416 364308 196504
rect 364416 196416 364596 196504
rect 364704 196416 364884 196504
rect 364992 196416 365172 196504
rect 365280 196416 365460 196504
rect 365714 196416 365894 196504
rect 366002 196416 366182 196504
rect 366290 196416 366470 196504
rect 366578 196416 366758 196504
rect 366866 196416 367046 196504
rect 367154 196416 367334 196504
rect 367442 196416 367622 196504
rect 367730 196416 367910 196504
rect 243214 196200 243394 196288
rect 243502 196200 243682 196288
rect 243790 196200 243970 196288
rect 244078 196200 244258 196288
rect 244366 196200 244546 196288
rect 244654 196200 244834 196288
rect 244942 196200 245122 196288
rect 245230 196200 245410 196288
rect 245664 196200 245844 196288
rect 245952 196200 246132 196288
rect 246240 196200 246420 196288
rect 246528 196200 246708 196288
rect 246816 196200 246996 196288
rect 247104 196200 247284 196288
rect 247392 196200 247572 196288
rect 247680 196200 247860 196288
rect 248114 196200 248294 196288
rect 248402 196200 248582 196288
rect 248690 196200 248870 196288
rect 248978 196200 249158 196288
rect 249266 196200 249446 196288
rect 249554 196200 249734 196288
rect 249842 196200 250022 196288
rect 250130 196200 250310 196288
rect 250564 196200 250744 196288
rect 360436 196200 360560 196288
rect 360814 196200 360994 196288
rect 361102 196200 361282 196288
rect 361390 196200 361570 196288
rect 361678 196200 361858 196288
rect 361966 196200 362146 196288
rect 362254 196200 362434 196288
rect 362542 196200 362722 196288
rect 362830 196200 363010 196288
rect 363264 196200 363444 196288
rect 363552 196200 363732 196288
rect 363840 196200 364020 196288
rect 364128 196200 364308 196288
rect 364416 196200 364596 196288
rect 364704 196200 364884 196288
rect 364992 196200 365172 196288
rect 365280 196200 365460 196288
rect 365714 196200 365894 196288
rect 366002 196200 366182 196288
rect 366290 196200 366470 196288
rect 366578 196200 366758 196288
rect 366866 196200 367046 196288
rect 367154 196200 367334 196288
rect 367442 196200 367622 196288
rect 367730 196200 367910 196288
rect 243214 195724 243394 195812
rect 243502 195724 243682 195812
rect 243790 195724 243970 195812
rect 244078 195724 244258 195812
rect 244366 195724 244546 195812
rect 244654 195724 244834 195812
rect 244942 195724 245122 195812
rect 245230 195724 245410 195812
rect 245664 195724 245844 195812
rect 245952 195724 246132 195812
rect 246240 195724 246420 195812
rect 246528 195724 246708 195812
rect 246816 195724 246996 195812
rect 247104 195724 247284 195812
rect 247392 195724 247572 195812
rect 247680 195724 247860 195812
rect 248114 195724 248294 195812
rect 248402 195724 248582 195812
rect 248690 195724 248870 195812
rect 248978 195724 249158 195812
rect 249266 195724 249446 195812
rect 249554 195724 249734 195812
rect 249842 195724 250022 195812
rect 250130 195724 250310 195812
rect 250564 195724 250744 195812
rect 360436 195724 360560 195812
rect 360814 195724 360994 195812
rect 361102 195724 361282 195812
rect 361390 195724 361570 195812
rect 361678 195724 361858 195812
rect 361966 195724 362146 195812
rect 362254 195724 362434 195812
rect 362542 195724 362722 195812
rect 362830 195724 363010 195812
rect 363264 195724 363444 195812
rect 363552 195724 363732 195812
rect 363840 195724 364020 195812
rect 364128 195724 364308 195812
rect 364416 195724 364596 195812
rect 364704 195724 364884 195812
rect 364992 195724 365172 195812
rect 365280 195724 365460 195812
rect 365714 195724 365894 195812
rect 366002 195724 366182 195812
rect 366290 195724 366470 195812
rect 366578 195724 366758 195812
rect 366866 195724 367046 195812
rect 367154 195724 367334 195812
rect 367442 195724 367622 195812
rect 367730 195724 367910 195812
rect 243214 195508 243394 195596
rect 243502 195508 243682 195596
rect 243790 195508 243970 195596
rect 244078 195508 244258 195596
rect 244366 195508 244546 195596
rect 244654 195508 244834 195596
rect 244942 195508 245122 195596
rect 245230 195508 245410 195596
rect 245664 195508 245844 195596
rect 245952 195508 246132 195596
rect 246240 195508 246420 195596
rect 246528 195508 246708 195596
rect 246816 195508 246996 195596
rect 247104 195508 247284 195596
rect 247392 195508 247572 195596
rect 247680 195508 247860 195596
rect 248114 195508 248294 195596
rect 248402 195508 248582 195596
rect 248690 195508 248870 195596
rect 248978 195508 249158 195596
rect 249266 195508 249446 195596
rect 249554 195508 249734 195596
rect 249842 195508 250022 195596
rect 250130 195508 250310 195596
rect 250564 195508 250744 195596
rect 360436 195508 360560 195596
rect 360814 195508 360994 195596
rect 361102 195508 361282 195596
rect 361390 195508 361570 195596
rect 361678 195508 361858 195596
rect 361966 195508 362146 195596
rect 362254 195508 362434 195596
rect 362542 195508 362722 195596
rect 362830 195508 363010 195596
rect 363264 195508 363444 195596
rect 363552 195508 363732 195596
rect 363840 195508 364020 195596
rect 364128 195508 364308 195596
rect 364416 195508 364596 195596
rect 364704 195508 364884 195596
rect 364992 195508 365172 195596
rect 365280 195508 365460 195596
rect 365714 195508 365894 195596
rect 366002 195508 366182 195596
rect 366290 195508 366470 195596
rect 366578 195508 366758 195596
rect 366866 195508 367046 195596
rect 367154 195508 367334 195596
rect 367442 195508 367622 195596
rect 367730 195508 367910 195596
rect 243214 195032 243394 195120
rect 243502 195032 243682 195120
rect 243790 195032 243970 195120
rect 244078 195032 244258 195120
rect 244366 195032 244546 195120
rect 244654 195032 244834 195120
rect 244942 195032 245122 195120
rect 245230 195032 245410 195120
rect 245664 195032 245844 195120
rect 245952 195032 246132 195120
rect 246240 195032 246420 195120
rect 246528 195032 246708 195120
rect 246816 195032 246996 195120
rect 247104 195032 247284 195120
rect 247392 195032 247572 195120
rect 247680 195032 247860 195120
rect 248114 195032 248294 195120
rect 248402 195032 248582 195120
rect 248690 195032 248870 195120
rect 248978 195032 249158 195120
rect 249266 195032 249446 195120
rect 249554 195032 249734 195120
rect 249842 195032 250022 195120
rect 250130 195032 250310 195120
rect 250564 195032 250744 195120
rect 360436 195032 360560 195120
rect 360814 195032 360994 195120
rect 361102 195032 361282 195120
rect 361390 195032 361570 195120
rect 361678 195032 361858 195120
rect 361966 195032 362146 195120
rect 362254 195032 362434 195120
rect 362542 195032 362722 195120
rect 362830 195032 363010 195120
rect 363264 195032 363444 195120
rect 363552 195032 363732 195120
rect 363840 195032 364020 195120
rect 364128 195032 364308 195120
rect 364416 195032 364596 195120
rect 364704 195032 364884 195120
rect 364992 195032 365172 195120
rect 365280 195032 365460 195120
rect 365714 195032 365894 195120
rect 366002 195032 366182 195120
rect 366290 195032 366470 195120
rect 366578 195032 366758 195120
rect 366866 195032 367046 195120
rect 367154 195032 367334 195120
rect 367442 195032 367622 195120
rect 367730 195032 367910 195120
rect 243214 194816 243394 194904
rect 243502 194816 243682 194904
rect 243790 194816 243970 194904
rect 244078 194816 244258 194904
rect 244366 194816 244546 194904
rect 244654 194816 244834 194904
rect 244942 194816 245122 194904
rect 245230 194816 245410 194904
rect 245664 194816 245844 194904
rect 245952 194816 246132 194904
rect 246240 194816 246420 194904
rect 246528 194816 246708 194904
rect 246816 194816 246996 194904
rect 247104 194816 247284 194904
rect 247392 194816 247572 194904
rect 247680 194816 247860 194904
rect 248114 194816 248294 194904
rect 248402 194816 248582 194904
rect 248690 194816 248870 194904
rect 248978 194816 249158 194904
rect 249266 194816 249446 194904
rect 249554 194816 249734 194904
rect 249842 194816 250022 194904
rect 250130 194816 250310 194904
rect 250564 194816 250744 194904
rect 360436 194816 360560 194904
rect 360814 194816 360994 194904
rect 361102 194816 361282 194904
rect 361390 194816 361570 194904
rect 361678 194816 361858 194904
rect 361966 194816 362146 194904
rect 362254 194816 362434 194904
rect 362542 194816 362722 194904
rect 362830 194816 363010 194904
rect 363264 194816 363444 194904
rect 363552 194816 363732 194904
rect 363840 194816 364020 194904
rect 364128 194816 364308 194904
rect 364416 194816 364596 194904
rect 364704 194816 364884 194904
rect 364992 194816 365172 194904
rect 365280 194816 365460 194904
rect 365714 194816 365894 194904
rect 366002 194816 366182 194904
rect 366290 194816 366470 194904
rect 366578 194816 366758 194904
rect 366866 194816 367046 194904
rect 367154 194816 367334 194904
rect 367442 194816 367622 194904
rect 367730 194816 367910 194904
rect 243214 194340 243394 194428
rect 243502 194340 243682 194428
rect 243790 194340 243970 194428
rect 244078 194340 244258 194428
rect 244366 194340 244546 194428
rect 244654 194340 244834 194428
rect 244942 194340 245122 194428
rect 245230 194340 245410 194428
rect 245664 194340 245844 194428
rect 245952 194340 246132 194428
rect 246240 194340 246420 194428
rect 246528 194340 246708 194428
rect 246816 194340 246996 194428
rect 247104 194340 247284 194428
rect 247392 194340 247572 194428
rect 247680 194340 247860 194428
rect 248114 194340 248294 194428
rect 248402 194340 248582 194428
rect 248690 194340 248870 194428
rect 248978 194340 249158 194428
rect 249266 194340 249446 194428
rect 249554 194340 249734 194428
rect 249842 194340 250022 194428
rect 250130 194340 250310 194428
rect 250564 194340 250744 194428
rect 360436 194340 360560 194428
rect 360814 194340 360994 194428
rect 361102 194340 361282 194428
rect 361390 194340 361570 194428
rect 361678 194340 361858 194428
rect 361966 194340 362146 194428
rect 362254 194340 362434 194428
rect 362542 194340 362722 194428
rect 362830 194340 363010 194428
rect 363264 194340 363444 194428
rect 363552 194340 363732 194428
rect 363840 194340 364020 194428
rect 364128 194340 364308 194428
rect 364416 194340 364596 194428
rect 364704 194340 364884 194428
rect 364992 194340 365172 194428
rect 365280 194340 365460 194428
rect 365714 194340 365894 194428
rect 366002 194340 366182 194428
rect 366290 194340 366470 194428
rect 366578 194340 366758 194428
rect 366866 194340 367046 194428
rect 367154 194340 367334 194428
rect 367442 194340 367622 194428
rect 367730 194340 367910 194428
rect 243214 193866 243394 193954
rect 243502 193866 243682 193954
rect 243790 193866 243970 193954
rect 244078 193866 244258 193954
rect 244366 193866 244546 193954
rect 244654 193866 244834 193954
rect 244942 193866 245122 193954
rect 245230 193866 245410 193954
rect 245664 193866 245844 193954
rect 245952 193866 246132 193954
rect 246240 193866 246420 193954
rect 246528 193866 246708 193954
rect 246816 193866 246996 193954
rect 247104 193866 247284 193954
rect 247392 193866 247572 193954
rect 247680 193866 247860 193954
rect 248114 193866 248294 193954
rect 248402 193866 248582 193954
rect 248690 193866 248870 193954
rect 248978 193866 249158 193954
rect 249266 193866 249446 193954
rect 249554 193866 249734 193954
rect 249842 193866 250022 193954
rect 250130 193866 250310 193954
rect 250564 193866 250744 193954
rect 360436 193866 360560 193954
rect 360814 193866 360994 193954
rect 361102 193866 361282 193954
rect 361390 193866 361570 193954
rect 361678 193866 361858 193954
rect 361966 193866 362146 193954
rect 362254 193866 362434 193954
rect 362542 193866 362722 193954
rect 362830 193866 363010 193954
rect 363264 193866 363444 193954
rect 363552 193866 363732 193954
rect 363840 193866 364020 193954
rect 364128 193866 364308 193954
rect 364416 193866 364596 193954
rect 364704 193866 364884 193954
rect 364992 193866 365172 193954
rect 365280 193866 365460 193954
rect 365714 193866 365894 193954
rect 366002 193866 366182 193954
rect 366290 193866 366470 193954
rect 366578 193866 366758 193954
rect 366866 193866 367046 193954
rect 367154 193866 367334 193954
rect 367442 193866 367622 193954
rect 367730 193866 367910 193954
rect 243214 193390 243394 193478
rect 243502 193390 243682 193478
rect 243790 193390 243970 193478
rect 244078 193390 244258 193478
rect 244366 193390 244546 193478
rect 244654 193390 244834 193478
rect 244942 193390 245122 193478
rect 245230 193390 245410 193478
rect 245664 193390 245844 193478
rect 245952 193390 246132 193478
rect 246240 193390 246420 193478
rect 246528 193390 246708 193478
rect 246816 193390 246996 193478
rect 247104 193390 247284 193478
rect 247392 193390 247572 193478
rect 247680 193390 247860 193478
rect 248114 193390 248294 193478
rect 248402 193390 248582 193478
rect 248690 193390 248870 193478
rect 248978 193390 249158 193478
rect 249266 193390 249446 193478
rect 249554 193390 249734 193478
rect 249842 193390 250022 193478
rect 250130 193390 250310 193478
rect 250564 193390 250744 193478
rect 360436 193390 360560 193478
rect 360814 193390 360994 193478
rect 361102 193390 361282 193478
rect 361390 193390 361570 193478
rect 361678 193390 361858 193478
rect 361966 193390 362146 193478
rect 362254 193390 362434 193478
rect 362542 193390 362722 193478
rect 362830 193390 363010 193478
rect 363264 193390 363444 193478
rect 363552 193390 363732 193478
rect 363840 193390 364020 193478
rect 364128 193390 364308 193478
rect 364416 193390 364596 193478
rect 364704 193390 364884 193478
rect 364992 193390 365172 193478
rect 365280 193390 365460 193478
rect 365714 193390 365894 193478
rect 366002 193390 366182 193478
rect 366290 193390 366470 193478
rect 366578 193390 366758 193478
rect 366866 193390 367046 193478
rect 367154 193390 367334 193478
rect 367442 193390 367622 193478
rect 367730 193390 367910 193478
rect 243214 193174 243394 193262
rect 243502 193174 243682 193262
rect 243790 193174 243970 193262
rect 244078 193174 244258 193262
rect 244366 193174 244546 193262
rect 244654 193174 244834 193262
rect 244942 193174 245122 193262
rect 245230 193174 245410 193262
rect 245664 193174 245844 193262
rect 245952 193174 246132 193262
rect 246240 193174 246420 193262
rect 246528 193174 246708 193262
rect 246816 193174 246996 193262
rect 247104 193174 247284 193262
rect 247392 193174 247572 193262
rect 247680 193174 247860 193262
rect 248114 193174 248294 193262
rect 248402 193174 248582 193262
rect 248690 193174 248870 193262
rect 248978 193174 249158 193262
rect 249266 193174 249446 193262
rect 249554 193174 249734 193262
rect 249842 193174 250022 193262
rect 250130 193174 250310 193262
rect 250564 193174 250744 193262
rect 360436 193174 360560 193262
rect 360814 193174 360994 193262
rect 361102 193174 361282 193262
rect 361390 193174 361570 193262
rect 361678 193174 361858 193262
rect 361966 193174 362146 193262
rect 362254 193174 362434 193262
rect 362542 193174 362722 193262
rect 362830 193174 363010 193262
rect 363264 193174 363444 193262
rect 363552 193174 363732 193262
rect 363840 193174 364020 193262
rect 364128 193174 364308 193262
rect 364416 193174 364596 193262
rect 364704 193174 364884 193262
rect 364992 193174 365172 193262
rect 365280 193174 365460 193262
rect 365714 193174 365894 193262
rect 366002 193174 366182 193262
rect 366290 193174 366470 193262
rect 366578 193174 366758 193262
rect 366866 193174 367046 193262
rect 367154 193174 367334 193262
rect 367442 193174 367622 193262
rect 367730 193174 367910 193262
rect 243214 192698 243394 192786
rect 243502 192698 243682 192786
rect 243790 192698 243970 192786
rect 244078 192698 244258 192786
rect 244366 192698 244546 192786
rect 244654 192698 244834 192786
rect 244942 192698 245122 192786
rect 245230 192698 245410 192786
rect 245664 192698 245844 192786
rect 245952 192698 246132 192786
rect 246240 192698 246420 192786
rect 246528 192698 246708 192786
rect 246816 192698 246996 192786
rect 247104 192698 247284 192786
rect 247392 192698 247572 192786
rect 247680 192698 247860 192786
rect 248114 192698 248294 192786
rect 248402 192698 248582 192786
rect 248690 192698 248870 192786
rect 248978 192698 249158 192786
rect 249266 192698 249446 192786
rect 249554 192698 249734 192786
rect 249842 192698 250022 192786
rect 250130 192698 250310 192786
rect 250564 192698 250744 192786
rect 360436 192698 360560 192786
rect 360814 192698 360994 192786
rect 361102 192698 361282 192786
rect 361390 192698 361570 192786
rect 361678 192698 361858 192786
rect 361966 192698 362146 192786
rect 362254 192698 362434 192786
rect 362542 192698 362722 192786
rect 362830 192698 363010 192786
rect 363264 192698 363444 192786
rect 363552 192698 363732 192786
rect 363840 192698 364020 192786
rect 364128 192698 364308 192786
rect 364416 192698 364596 192786
rect 364704 192698 364884 192786
rect 364992 192698 365172 192786
rect 365280 192698 365460 192786
rect 365714 192698 365894 192786
rect 366002 192698 366182 192786
rect 366290 192698 366470 192786
rect 366578 192698 366758 192786
rect 366866 192698 367046 192786
rect 367154 192698 367334 192786
rect 367442 192698 367622 192786
rect 367730 192698 367910 192786
rect 243214 192482 243394 192570
rect 243502 192482 243682 192570
rect 243790 192482 243970 192570
rect 244078 192482 244258 192570
rect 244366 192482 244546 192570
rect 244654 192482 244834 192570
rect 244942 192482 245122 192570
rect 245230 192482 245410 192570
rect 245664 192482 245844 192570
rect 245952 192482 246132 192570
rect 246240 192482 246420 192570
rect 246528 192482 246708 192570
rect 246816 192482 246996 192570
rect 247104 192482 247284 192570
rect 247392 192482 247572 192570
rect 247680 192482 247860 192570
rect 248114 192482 248294 192570
rect 248402 192482 248582 192570
rect 248690 192482 248870 192570
rect 248978 192482 249158 192570
rect 249266 192482 249446 192570
rect 249554 192482 249734 192570
rect 249842 192482 250022 192570
rect 250130 192482 250310 192570
rect 250564 192482 250744 192570
rect 360436 192482 360560 192570
rect 360814 192482 360994 192570
rect 361102 192482 361282 192570
rect 361390 192482 361570 192570
rect 361678 192482 361858 192570
rect 361966 192482 362146 192570
rect 362254 192482 362434 192570
rect 362542 192482 362722 192570
rect 362830 192482 363010 192570
rect 363264 192482 363444 192570
rect 363552 192482 363732 192570
rect 363840 192482 364020 192570
rect 364128 192482 364308 192570
rect 364416 192482 364596 192570
rect 364704 192482 364884 192570
rect 364992 192482 365172 192570
rect 365280 192482 365460 192570
rect 365714 192482 365894 192570
rect 366002 192482 366182 192570
rect 366290 192482 366470 192570
rect 366578 192482 366758 192570
rect 366866 192482 367046 192570
rect 367154 192482 367334 192570
rect 367442 192482 367622 192570
rect 367730 192482 367910 192570
rect 243214 192006 243394 192094
rect 243502 192006 243682 192094
rect 243790 192006 243970 192094
rect 244078 192006 244258 192094
rect 244366 192006 244546 192094
rect 244654 192006 244834 192094
rect 244942 192006 245122 192094
rect 245230 192006 245410 192094
rect 245664 192006 245844 192094
rect 245952 192006 246132 192094
rect 246240 192006 246420 192094
rect 246528 192006 246708 192094
rect 246816 192006 246996 192094
rect 247104 192006 247284 192094
rect 247392 192006 247572 192094
rect 247680 192006 247860 192094
rect 248114 192006 248294 192094
rect 248402 192006 248582 192094
rect 248690 192006 248870 192094
rect 248978 192006 249158 192094
rect 249266 192006 249446 192094
rect 249554 192006 249734 192094
rect 249842 192006 250022 192094
rect 250130 192006 250310 192094
rect 250564 192006 250744 192094
rect 360436 192006 360560 192094
rect 360814 192006 360994 192094
rect 361102 192006 361282 192094
rect 361390 192006 361570 192094
rect 361678 192006 361858 192094
rect 361966 192006 362146 192094
rect 362254 192006 362434 192094
rect 362542 192006 362722 192094
rect 362830 192006 363010 192094
rect 363264 192006 363444 192094
rect 363552 192006 363732 192094
rect 363840 192006 364020 192094
rect 364128 192006 364308 192094
rect 364416 192006 364596 192094
rect 364704 192006 364884 192094
rect 364992 192006 365172 192094
rect 365280 192006 365460 192094
rect 365714 192006 365894 192094
rect 366002 192006 366182 192094
rect 366290 192006 366470 192094
rect 366578 192006 366758 192094
rect 366866 192006 367046 192094
rect 367154 192006 367334 192094
rect 367442 192006 367622 192094
rect 367730 192006 367910 192094
rect 243214 191790 243394 191878
rect 243502 191790 243682 191878
rect 243790 191790 243970 191878
rect 244078 191790 244258 191878
rect 244366 191790 244546 191878
rect 244654 191790 244834 191878
rect 244942 191790 245122 191878
rect 245230 191790 245410 191878
rect 245664 191790 245844 191878
rect 245952 191790 246132 191878
rect 246240 191790 246420 191878
rect 246528 191790 246708 191878
rect 246816 191790 246996 191878
rect 247104 191790 247284 191878
rect 247392 191790 247572 191878
rect 247680 191790 247860 191878
rect 248114 191790 248294 191878
rect 248402 191790 248582 191878
rect 248690 191790 248870 191878
rect 248978 191790 249158 191878
rect 249266 191790 249446 191878
rect 249554 191790 249734 191878
rect 249842 191790 250022 191878
rect 250130 191790 250310 191878
rect 250564 191790 250744 191878
rect 360436 191790 360560 191878
rect 360814 191790 360994 191878
rect 361102 191790 361282 191878
rect 361390 191790 361570 191878
rect 361678 191790 361858 191878
rect 361966 191790 362146 191878
rect 362254 191790 362434 191878
rect 362542 191790 362722 191878
rect 362830 191790 363010 191878
rect 363264 191790 363444 191878
rect 363552 191790 363732 191878
rect 363840 191790 364020 191878
rect 364128 191790 364308 191878
rect 364416 191790 364596 191878
rect 364704 191790 364884 191878
rect 364992 191790 365172 191878
rect 365280 191790 365460 191878
rect 365714 191790 365894 191878
rect 366002 191790 366182 191878
rect 366290 191790 366470 191878
rect 366578 191790 366758 191878
rect 366866 191790 367046 191878
rect 367154 191790 367334 191878
rect 367442 191790 367622 191878
rect 367730 191790 367910 191878
rect 243214 191314 243394 191402
rect 243502 191314 243682 191402
rect 243790 191314 243970 191402
rect 244078 191314 244258 191402
rect 244366 191314 244546 191402
rect 244654 191314 244834 191402
rect 244942 191314 245122 191402
rect 245230 191314 245410 191402
rect 245664 191314 245844 191402
rect 245952 191314 246132 191402
rect 246240 191314 246420 191402
rect 246528 191314 246708 191402
rect 246816 191314 246996 191402
rect 247104 191314 247284 191402
rect 247392 191314 247572 191402
rect 247680 191314 247860 191402
rect 248114 191314 248294 191402
rect 248402 191314 248582 191402
rect 248690 191314 248870 191402
rect 248978 191314 249158 191402
rect 249266 191314 249446 191402
rect 249554 191314 249734 191402
rect 249842 191314 250022 191402
rect 250130 191314 250310 191402
rect 250564 191314 250744 191402
rect 360436 191314 360560 191402
rect 360814 191314 360994 191402
rect 361102 191314 361282 191402
rect 361390 191314 361570 191402
rect 361678 191314 361858 191402
rect 361966 191314 362146 191402
rect 362254 191314 362434 191402
rect 362542 191314 362722 191402
rect 362830 191314 363010 191402
rect 363264 191314 363444 191402
rect 363552 191314 363732 191402
rect 363840 191314 364020 191402
rect 364128 191314 364308 191402
rect 364416 191314 364596 191402
rect 364704 191314 364884 191402
rect 364992 191314 365172 191402
rect 365280 191314 365460 191402
rect 365714 191314 365894 191402
rect 366002 191314 366182 191402
rect 366290 191314 366470 191402
rect 366578 191314 366758 191402
rect 366866 191314 367046 191402
rect 367154 191314 367334 191402
rect 367442 191314 367622 191402
rect 367730 191314 367910 191402
rect 243214 190840 243394 190928
rect 243502 190840 243682 190928
rect 243790 190840 243970 190928
rect 244078 190840 244258 190928
rect 244366 190840 244546 190928
rect 244654 190840 244834 190928
rect 244942 190840 245122 190928
rect 245230 190840 245410 190928
rect 245664 190840 245844 190928
rect 245952 190840 246132 190928
rect 246240 190840 246420 190928
rect 246528 190840 246708 190928
rect 246816 190840 246996 190928
rect 247104 190840 247284 190928
rect 247392 190840 247572 190928
rect 247680 190840 247860 190928
rect 248114 190840 248294 190928
rect 248402 190840 248582 190928
rect 248690 190840 248870 190928
rect 248978 190840 249158 190928
rect 249266 190840 249446 190928
rect 249554 190840 249734 190928
rect 249842 190840 250022 190928
rect 250130 190840 250310 190928
rect 250564 190840 250744 190928
rect 360436 190840 360560 190928
rect 360814 190840 360994 190928
rect 361102 190840 361282 190928
rect 361390 190840 361570 190928
rect 361678 190840 361858 190928
rect 361966 190840 362146 190928
rect 362254 190840 362434 190928
rect 362542 190840 362722 190928
rect 362830 190840 363010 190928
rect 363264 190840 363444 190928
rect 363552 190840 363732 190928
rect 363840 190840 364020 190928
rect 364128 190840 364308 190928
rect 364416 190840 364596 190928
rect 364704 190840 364884 190928
rect 364992 190840 365172 190928
rect 365280 190840 365460 190928
rect 365714 190840 365894 190928
rect 366002 190840 366182 190928
rect 366290 190840 366470 190928
rect 366578 190840 366758 190928
rect 366866 190840 367046 190928
rect 367154 190840 367334 190928
rect 367442 190840 367622 190928
rect 367730 190840 367910 190928
rect 243214 190364 243394 190452
rect 243502 190364 243682 190452
rect 243790 190364 243970 190452
rect 244078 190364 244258 190452
rect 244366 190364 244546 190452
rect 244654 190364 244834 190452
rect 244942 190364 245122 190452
rect 245230 190364 245410 190452
rect 245664 190364 245844 190452
rect 245952 190364 246132 190452
rect 246240 190364 246420 190452
rect 246528 190364 246708 190452
rect 246816 190364 246996 190452
rect 247104 190364 247284 190452
rect 247392 190364 247572 190452
rect 247680 190364 247860 190452
rect 248114 190364 248294 190452
rect 248402 190364 248582 190452
rect 248690 190364 248870 190452
rect 248978 190364 249158 190452
rect 249266 190364 249446 190452
rect 249554 190364 249734 190452
rect 249842 190364 250022 190452
rect 250130 190364 250310 190452
rect 250564 190364 250744 190452
rect 360436 190364 360560 190452
rect 360814 190364 360994 190452
rect 361102 190364 361282 190452
rect 361390 190364 361570 190452
rect 361678 190364 361858 190452
rect 361966 190364 362146 190452
rect 362254 190364 362434 190452
rect 362542 190364 362722 190452
rect 362830 190364 363010 190452
rect 363264 190364 363444 190452
rect 363552 190364 363732 190452
rect 363840 190364 364020 190452
rect 364128 190364 364308 190452
rect 364416 190364 364596 190452
rect 364704 190364 364884 190452
rect 364992 190364 365172 190452
rect 365280 190364 365460 190452
rect 365714 190364 365894 190452
rect 366002 190364 366182 190452
rect 366290 190364 366470 190452
rect 366578 190364 366758 190452
rect 366866 190364 367046 190452
rect 367154 190364 367334 190452
rect 367442 190364 367622 190452
rect 367730 190364 367910 190452
rect 243214 190148 243394 190236
rect 243502 190148 243682 190236
rect 243790 190148 243970 190236
rect 244078 190148 244258 190236
rect 244366 190148 244546 190236
rect 244654 190148 244834 190236
rect 244942 190148 245122 190236
rect 245230 190148 245410 190236
rect 245664 190148 245844 190236
rect 245952 190148 246132 190236
rect 246240 190148 246420 190236
rect 246528 190148 246708 190236
rect 246816 190148 246996 190236
rect 247104 190148 247284 190236
rect 247392 190148 247572 190236
rect 247680 190148 247860 190236
rect 248114 190148 248294 190236
rect 248402 190148 248582 190236
rect 248690 190148 248870 190236
rect 248978 190148 249158 190236
rect 249266 190148 249446 190236
rect 249554 190148 249734 190236
rect 249842 190148 250022 190236
rect 250130 190148 250310 190236
rect 250564 190148 250744 190236
rect 360436 190148 360560 190236
rect 360814 190148 360994 190236
rect 361102 190148 361282 190236
rect 361390 190148 361570 190236
rect 361678 190148 361858 190236
rect 361966 190148 362146 190236
rect 362254 190148 362434 190236
rect 362542 190148 362722 190236
rect 362830 190148 363010 190236
rect 363264 190148 363444 190236
rect 363552 190148 363732 190236
rect 363840 190148 364020 190236
rect 364128 190148 364308 190236
rect 364416 190148 364596 190236
rect 364704 190148 364884 190236
rect 364992 190148 365172 190236
rect 365280 190148 365460 190236
rect 365714 190148 365894 190236
rect 366002 190148 366182 190236
rect 366290 190148 366470 190236
rect 366578 190148 366758 190236
rect 366866 190148 367046 190236
rect 367154 190148 367334 190236
rect 367442 190148 367622 190236
rect 367730 190148 367910 190236
rect 243214 189672 243394 189760
rect 243502 189672 243682 189760
rect 243790 189672 243970 189760
rect 244078 189672 244258 189760
rect 244366 189672 244546 189760
rect 244654 189672 244834 189760
rect 244942 189672 245122 189760
rect 245230 189672 245410 189760
rect 245664 189672 245844 189760
rect 245952 189672 246132 189760
rect 246240 189672 246420 189760
rect 246528 189672 246708 189760
rect 246816 189672 246996 189760
rect 247104 189672 247284 189760
rect 247392 189672 247572 189760
rect 247680 189672 247860 189760
rect 248114 189672 248294 189760
rect 248402 189672 248582 189760
rect 248690 189672 248870 189760
rect 248978 189672 249158 189760
rect 249266 189672 249446 189760
rect 249554 189672 249734 189760
rect 249842 189672 250022 189760
rect 250130 189672 250310 189760
rect 250564 189672 250744 189760
rect 360436 189672 360560 189760
rect 360814 189672 360994 189760
rect 361102 189672 361282 189760
rect 361390 189672 361570 189760
rect 361678 189672 361858 189760
rect 361966 189672 362146 189760
rect 362254 189672 362434 189760
rect 362542 189672 362722 189760
rect 362830 189672 363010 189760
rect 363264 189672 363444 189760
rect 363552 189672 363732 189760
rect 363840 189672 364020 189760
rect 364128 189672 364308 189760
rect 364416 189672 364596 189760
rect 364704 189672 364884 189760
rect 364992 189672 365172 189760
rect 365280 189672 365460 189760
rect 365714 189672 365894 189760
rect 366002 189672 366182 189760
rect 366290 189672 366470 189760
rect 366578 189672 366758 189760
rect 366866 189672 367046 189760
rect 367154 189672 367334 189760
rect 367442 189672 367622 189760
rect 367730 189672 367910 189760
rect 243214 189456 243394 189544
rect 243502 189456 243682 189544
rect 243790 189456 243970 189544
rect 244078 189456 244258 189544
rect 244366 189456 244546 189544
rect 244654 189456 244834 189544
rect 244942 189456 245122 189544
rect 245230 189456 245410 189544
rect 245664 189456 245844 189544
rect 245952 189456 246132 189544
rect 246240 189456 246420 189544
rect 246528 189456 246708 189544
rect 246816 189456 246996 189544
rect 247104 189456 247284 189544
rect 247392 189456 247572 189544
rect 247680 189456 247860 189544
rect 248114 189456 248294 189544
rect 248402 189456 248582 189544
rect 248690 189456 248870 189544
rect 248978 189456 249158 189544
rect 249266 189456 249446 189544
rect 249554 189456 249734 189544
rect 249842 189456 250022 189544
rect 250130 189456 250310 189544
rect 250564 189456 250744 189544
rect 360436 189456 360560 189544
rect 360814 189456 360994 189544
rect 361102 189456 361282 189544
rect 361390 189456 361570 189544
rect 361678 189456 361858 189544
rect 361966 189456 362146 189544
rect 362254 189456 362434 189544
rect 362542 189456 362722 189544
rect 362830 189456 363010 189544
rect 363264 189456 363444 189544
rect 363552 189456 363732 189544
rect 363840 189456 364020 189544
rect 364128 189456 364308 189544
rect 364416 189456 364596 189544
rect 364704 189456 364884 189544
rect 364992 189456 365172 189544
rect 365280 189456 365460 189544
rect 365714 189456 365894 189544
rect 366002 189456 366182 189544
rect 366290 189456 366470 189544
rect 366578 189456 366758 189544
rect 366866 189456 367046 189544
rect 367154 189456 367334 189544
rect 367442 189456 367622 189544
rect 367730 189456 367910 189544
rect 243214 188980 243394 189068
rect 243502 188980 243682 189068
rect 243790 188980 243970 189068
rect 244078 188980 244258 189068
rect 244366 188980 244546 189068
rect 244654 188980 244834 189068
rect 244942 188980 245122 189068
rect 245230 188980 245410 189068
rect 245664 188980 245844 189068
rect 245952 188980 246132 189068
rect 246240 188980 246420 189068
rect 246528 188980 246708 189068
rect 246816 188980 246996 189068
rect 247104 188980 247284 189068
rect 247392 188980 247572 189068
rect 247680 188980 247860 189068
rect 248114 188980 248294 189068
rect 248402 188980 248582 189068
rect 248690 188980 248870 189068
rect 248978 188980 249158 189068
rect 249266 188980 249446 189068
rect 249554 188980 249734 189068
rect 249842 188980 250022 189068
rect 250130 188980 250310 189068
rect 250564 188980 250744 189068
rect 360436 188980 360560 189068
rect 360814 188980 360994 189068
rect 361102 188980 361282 189068
rect 361390 188980 361570 189068
rect 361678 188980 361858 189068
rect 361966 188980 362146 189068
rect 362254 188980 362434 189068
rect 362542 188980 362722 189068
rect 362830 188980 363010 189068
rect 363264 188980 363444 189068
rect 363552 188980 363732 189068
rect 363840 188980 364020 189068
rect 364128 188980 364308 189068
rect 364416 188980 364596 189068
rect 364704 188980 364884 189068
rect 364992 188980 365172 189068
rect 365280 188980 365460 189068
rect 365714 188980 365894 189068
rect 366002 188980 366182 189068
rect 366290 188980 366470 189068
rect 366578 188980 366758 189068
rect 366866 188980 367046 189068
rect 367154 188980 367334 189068
rect 367442 188980 367622 189068
rect 367730 188980 367910 189068
rect 243214 188764 243394 188852
rect 243502 188764 243682 188852
rect 243790 188764 243970 188852
rect 244078 188764 244258 188852
rect 244366 188764 244546 188852
rect 244654 188764 244834 188852
rect 244942 188764 245122 188852
rect 245230 188764 245410 188852
rect 245664 188764 245844 188852
rect 245952 188764 246132 188852
rect 246240 188764 246420 188852
rect 246528 188764 246708 188852
rect 246816 188764 246996 188852
rect 247104 188764 247284 188852
rect 247392 188764 247572 188852
rect 247680 188764 247860 188852
rect 248114 188764 248294 188852
rect 248402 188764 248582 188852
rect 248690 188764 248870 188852
rect 248978 188764 249158 188852
rect 249266 188764 249446 188852
rect 249554 188764 249734 188852
rect 249842 188764 250022 188852
rect 250130 188764 250310 188852
rect 250564 188764 250744 188852
rect 360436 188764 360560 188852
rect 360814 188764 360994 188852
rect 361102 188764 361282 188852
rect 361390 188764 361570 188852
rect 361678 188764 361858 188852
rect 361966 188764 362146 188852
rect 362254 188764 362434 188852
rect 362542 188764 362722 188852
rect 362830 188764 363010 188852
rect 363264 188764 363444 188852
rect 363552 188764 363732 188852
rect 363840 188764 364020 188852
rect 364128 188764 364308 188852
rect 364416 188764 364596 188852
rect 364704 188764 364884 188852
rect 364992 188764 365172 188852
rect 365280 188764 365460 188852
rect 365714 188764 365894 188852
rect 366002 188764 366182 188852
rect 366290 188764 366470 188852
rect 366578 188764 366758 188852
rect 366866 188764 367046 188852
rect 367154 188764 367334 188852
rect 367442 188764 367622 188852
rect 367730 188764 367910 188852
rect 243214 188288 243394 188376
rect 243502 188288 243682 188376
rect 243790 188288 243970 188376
rect 244078 188288 244258 188376
rect 244366 188288 244546 188376
rect 244654 188288 244834 188376
rect 244942 188288 245122 188376
rect 245230 188288 245410 188376
rect 245664 188288 245844 188376
rect 245952 188288 246132 188376
rect 246240 188288 246420 188376
rect 246528 188288 246708 188376
rect 246816 188288 246996 188376
rect 247104 188288 247284 188376
rect 247392 188288 247572 188376
rect 247680 188288 247860 188376
rect 248114 188288 248294 188376
rect 248402 188288 248582 188376
rect 248690 188288 248870 188376
rect 248978 188288 249158 188376
rect 249266 188288 249446 188376
rect 249554 188288 249734 188376
rect 249842 188288 250022 188376
rect 250130 188288 250310 188376
rect 250564 188288 250744 188376
rect 360436 188288 360560 188376
rect 360814 188288 360994 188376
rect 361102 188288 361282 188376
rect 361390 188288 361570 188376
rect 361678 188288 361858 188376
rect 361966 188288 362146 188376
rect 362254 188288 362434 188376
rect 362542 188288 362722 188376
rect 362830 188288 363010 188376
rect 363264 188288 363444 188376
rect 363552 188288 363732 188376
rect 363840 188288 364020 188376
rect 364128 188288 364308 188376
rect 364416 188288 364596 188376
rect 364704 188288 364884 188376
rect 364992 188288 365172 188376
rect 365280 188288 365460 188376
rect 365714 188288 365894 188376
rect 366002 188288 366182 188376
rect 366290 188288 366470 188376
rect 366578 188288 366758 188376
rect 366866 188288 367046 188376
rect 367154 188288 367334 188376
rect 367442 188288 367622 188376
rect 367730 188288 367910 188376
rect 243214 187814 243394 187902
rect 243502 187814 243682 187902
rect 243790 187814 243970 187902
rect 244078 187814 244258 187902
rect 244366 187814 244546 187902
rect 244654 187814 244834 187902
rect 244942 187814 245122 187902
rect 245230 187814 245410 187902
rect 245664 187814 245844 187902
rect 245952 187814 246132 187902
rect 246240 187814 246420 187902
rect 246528 187814 246708 187902
rect 246816 187814 246996 187902
rect 247104 187814 247284 187902
rect 247392 187814 247572 187902
rect 247680 187814 247860 187902
rect 248114 187814 248294 187902
rect 248402 187814 248582 187902
rect 248690 187814 248870 187902
rect 248978 187814 249158 187902
rect 249266 187814 249446 187902
rect 249554 187814 249734 187902
rect 249842 187814 250022 187902
rect 250130 187814 250310 187902
rect 250564 187814 250744 187902
rect 360436 187814 360560 187902
rect 360814 187814 360994 187902
rect 361102 187814 361282 187902
rect 361390 187814 361570 187902
rect 361678 187814 361858 187902
rect 361966 187814 362146 187902
rect 362254 187814 362434 187902
rect 362542 187814 362722 187902
rect 362830 187814 363010 187902
rect 363264 187814 363444 187902
rect 363552 187814 363732 187902
rect 363840 187814 364020 187902
rect 364128 187814 364308 187902
rect 364416 187814 364596 187902
rect 364704 187814 364884 187902
rect 364992 187814 365172 187902
rect 365280 187814 365460 187902
rect 365714 187814 365894 187902
rect 366002 187814 366182 187902
rect 366290 187814 366470 187902
rect 366578 187814 366758 187902
rect 366866 187814 367046 187902
rect 367154 187814 367334 187902
rect 367442 187814 367622 187902
rect 367730 187814 367910 187902
rect 243214 187338 243394 187426
rect 243502 187338 243682 187426
rect 243790 187338 243970 187426
rect 244078 187338 244258 187426
rect 244366 187338 244546 187426
rect 244654 187338 244834 187426
rect 244942 187338 245122 187426
rect 245230 187338 245410 187426
rect 245664 187338 245844 187426
rect 245952 187338 246132 187426
rect 246240 187338 246420 187426
rect 246528 187338 246708 187426
rect 246816 187338 246996 187426
rect 247104 187338 247284 187426
rect 247392 187338 247572 187426
rect 247680 187338 247860 187426
rect 248114 187338 248294 187426
rect 248402 187338 248582 187426
rect 248690 187338 248870 187426
rect 248978 187338 249158 187426
rect 249266 187338 249446 187426
rect 249554 187338 249734 187426
rect 249842 187338 250022 187426
rect 250130 187338 250310 187426
rect 250564 187338 250744 187426
rect 360436 187338 360560 187426
rect 360814 187338 360994 187426
rect 361102 187338 361282 187426
rect 361390 187338 361570 187426
rect 361678 187338 361858 187426
rect 361966 187338 362146 187426
rect 362254 187338 362434 187426
rect 362542 187338 362722 187426
rect 362830 187338 363010 187426
rect 363264 187338 363444 187426
rect 363552 187338 363732 187426
rect 363840 187338 364020 187426
rect 364128 187338 364308 187426
rect 364416 187338 364596 187426
rect 364704 187338 364884 187426
rect 364992 187338 365172 187426
rect 365280 187338 365460 187426
rect 365714 187338 365894 187426
rect 366002 187338 366182 187426
rect 366290 187338 366470 187426
rect 366578 187338 366758 187426
rect 366866 187338 367046 187426
rect 367154 187338 367334 187426
rect 367442 187338 367622 187426
rect 367730 187338 367910 187426
rect 243214 187122 243394 187210
rect 243502 187122 243682 187210
rect 243790 187122 243970 187210
rect 244078 187122 244258 187210
rect 244366 187122 244546 187210
rect 244654 187122 244834 187210
rect 244942 187122 245122 187210
rect 245230 187122 245410 187210
rect 245664 187122 245844 187210
rect 245952 187122 246132 187210
rect 246240 187122 246420 187210
rect 246528 187122 246708 187210
rect 246816 187122 246996 187210
rect 247104 187122 247284 187210
rect 247392 187122 247572 187210
rect 247680 187122 247860 187210
rect 248114 187122 248294 187210
rect 248402 187122 248582 187210
rect 248690 187122 248870 187210
rect 248978 187122 249158 187210
rect 249266 187122 249446 187210
rect 249554 187122 249734 187210
rect 249842 187122 250022 187210
rect 250130 187122 250310 187210
rect 250564 187122 250744 187210
rect 360436 187122 360560 187210
rect 360814 187122 360994 187210
rect 361102 187122 361282 187210
rect 361390 187122 361570 187210
rect 361678 187122 361858 187210
rect 361966 187122 362146 187210
rect 362254 187122 362434 187210
rect 362542 187122 362722 187210
rect 362830 187122 363010 187210
rect 363264 187122 363444 187210
rect 363552 187122 363732 187210
rect 363840 187122 364020 187210
rect 364128 187122 364308 187210
rect 364416 187122 364596 187210
rect 364704 187122 364884 187210
rect 364992 187122 365172 187210
rect 365280 187122 365460 187210
rect 365714 187122 365894 187210
rect 366002 187122 366182 187210
rect 366290 187122 366470 187210
rect 366578 187122 366758 187210
rect 366866 187122 367046 187210
rect 367154 187122 367334 187210
rect 367442 187122 367622 187210
rect 367730 187122 367910 187210
rect 243214 186646 243394 186734
rect 243502 186646 243682 186734
rect 243790 186646 243970 186734
rect 244078 186646 244258 186734
rect 244366 186646 244546 186734
rect 244654 186646 244834 186734
rect 244942 186646 245122 186734
rect 245230 186646 245410 186734
rect 245664 186646 245844 186734
rect 245952 186646 246132 186734
rect 246240 186646 246420 186734
rect 246528 186646 246708 186734
rect 246816 186646 246996 186734
rect 247104 186646 247284 186734
rect 247392 186646 247572 186734
rect 247680 186646 247860 186734
rect 248114 186646 248294 186734
rect 248402 186646 248582 186734
rect 248690 186646 248870 186734
rect 248978 186646 249158 186734
rect 249266 186646 249446 186734
rect 249554 186646 249734 186734
rect 249842 186646 250022 186734
rect 250130 186646 250310 186734
rect 250564 186646 250744 186734
rect 360436 186646 360560 186734
rect 360814 186646 360994 186734
rect 361102 186646 361282 186734
rect 361390 186646 361570 186734
rect 361678 186646 361858 186734
rect 361966 186646 362146 186734
rect 362254 186646 362434 186734
rect 362542 186646 362722 186734
rect 362830 186646 363010 186734
rect 363264 186646 363444 186734
rect 363552 186646 363732 186734
rect 363840 186646 364020 186734
rect 364128 186646 364308 186734
rect 364416 186646 364596 186734
rect 364704 186646 364884 186734
rect 364992 186646 365172 186734
rect 365280 186646 365460 186734
rect 365714 186646 365894 186734
rect 366002 186646 366182 186734
rect 366290 186646 366470 186734
rect 366578 186646 366758 186734
rect 366866 186646 367046 186734
rect 367154 186646 367334 186734
rect 367442 186646 367622 186734
rect 367730 186646 367910 186734
rect 243214 186430 243394 186518
rect 243502 186430 243682 186518
rect 243790 186430 243970 186518
rect 244078 186430 244258 186518
rect 244366 186430 244546 186518
rect 244654 186430 244834 186518
rect 244942 186430 245122 186518
rect 245230 186430 245410 186518
rect 245664 186430 245844 186518
rect 245952 186430 246132 186518
rect 246240 186430 246420 186518
rect 246528 186430 246708 186518
rect 246816 186430 246996 186518
rect 247104 186430 247284 186518
rect 247392 186430 247572 186518
rect 247680 186430 247860 186518
rect 248114 186430 248294 186518
rect 248402 186430 248582 186518
rect 248690 186430 248870 186518
rect 248978 186430 249158 186518
rect 249266 186430 249446 186518
rect 249554 186430 249734 186518
rect 249842 186430 250022 186518
rect 250130 186430 250310 186518
rect 250564 186430 250744 186518
rect 360436 186430 360560 186518
rect 360814 186430 360994 186518
rect 361102 186430 361282 186518
rect 361390 186430 361570 186518
rect 361678 186430 361858 186518
rect 361966 186430 362146 186518
rect 362254 186430 362434 186518
rect 362542 186430 362722 186518
rect 362830 186430 363010 186518
rect 363264 186430 363444 186518
rect 363552 186430 363732 186518
rect 363840 186430 364020 186518
rect 364128 186430 364308 186518
rect 364416 186430 364596 186518
rect 364704 186430 364884 186518
rect 364992 186430 365172 186518
rect 365280 186430 365460 186518
rect 365714 186430 365894 186518
rect 366002 186430 366182 186518
rect 366290 186430 366470 186518
rect 366578 186430 366758 186518
rect 366866 186430 367046 186518
rect 367154 186430 367334 186518
rect 367442 186430 367622 186518
rect 367730 186430 367910 186518
rect 243214 185954 243394 186042
rect 243502 185954 243682 186042
rect 243790 185954 243970 186042
rect 244078 185954 244258 186042
rect 244366 185954 244546 186042
rect 244654 185954 244834 186042
rect 244942 185954 245122 186042
rect 245230 185954 245410 186042
rect 245664 185954 245844 186042
rect 245952 185954 246132 186042
rect 246240 185954 246420 186042
rect 246528 185954 246708 186042
rect 246816 185954 246996 186042
rect 247104 185954 247284 186042
rect 247392 185954 247572 186042
rect 247680 185954 247860 186042
rect 248114 185954 248294 186042
rect 248402 185954 248582 186042
rect 248690 185954 248870 186042
rect 248978 185954 249158 186042
rect 249266 185954 249446 186042
rect 249554 185954 249734 186042
rect 249842 185954 250022 186042
rect 250130 185954 250310 186042
rect 250564 185954 250744 186042
rect 360436 185954 360560 186042
rect 360814 185954 360994 186042
rect 361102 185954 361282 186042
rect 361390 185954 361570 186042
rect 361678 185954 361858 186042
rect 361966 185954 362146 186042
rect 362254 185954 362434 186042
rect 362542 185954 362722 186042
rect 362830 185954 363010 186042
rect 363264 185954 363444 186042
rect 363552 185954 363732 186042
rect 363840 185954 364020 186042
rect 364128 185954 364308 186042
rect 364416 185954 364596 186042
rect 364704 185954 364884 186042
rect 364992 185954 365172 186042
rect 365280 185954 365460 186042
rect 365714 185954 365894 186042
rect 366002 185954 366182 186042
rect 366290 185954 366470 186042
rect 366578 185954 366758 186042
rect 366866 185954 367046 186042
rect 367154 185954 367334 186042
rect 367442 185954 367622 186042
rect 367730 185954 367910 186042
rect 243214 185738 243394 185826
rect 243502 185738 243682 185826
rect 243790 185738 243970 185826
rect 244078 185738 244258 185826
rect 244366 185738 244546 185826
rect 244654 185738 244834 185826
rect 244942 185738 245122 185826
rect 245230 185738 245410 185826
rect 245664 185738 245844 185826
rect 245952 185738 246132 185826
rect 246240 185738 246420 185826
rect 246528 185738 246708 185826
rect 246816 185738 246996 185826
rect 247104 185738 247284 185826
rect 247392 185738 247572 185826
rect 247680 185738 247860 185826
rect 248114 185738 248294 185826
rect 248402 185738 248582 185826
rect 248690 185738 248870 185826
rect 248978 185738 249158 185826
rect 249266 185738 249446 185826
rect 249554 185738 249734 185826
rect 249842 185738 250022 185826
rect 250130 185738 250310 185826
rect 250564 185738 250744 185826
rect 360436 185738 360560 185826
rect 360814 185738 360994 185826
rect 361102 185738 361282 185826
rect 361390 185738 361570 185826
rect 361678 185738 361858 185826
rect 361966 185738 362146 185826
rect 362254 185738 362434 185826
rect 362542 185738 362722 185826
rect 362830 185738 363010 185826
rect 363264 185738 363444 185826
rect 363552 185738 363732 185826
rect 363840 185738 364020 185826
rect 364128 185738 364308 185826
rect 364416 185738 364596 185826
rect 364704 185738 364884 185826
rect 364992 185738 365172 185826
rect 365280 185738 365460 185826
rect 365714 185738 365894 185826
rect 366002 185738 366182 185826
rect 366290 185738 366470 185826
rect 366578 185738 366758 185826
rect 366866 185738 367046 185826
rect 367154 185738 367334 185826
rect 367442 185738 367622 185826
rect 367730 185738 367910 185826
rect 243214 185262 243394 185350
rect 243502 185262 243682 185350
rect 243790 185262 243970 185350
rect 244078 185262 244258 185350
rect 244366 185262 244546 185350
rect 244654 185262 244834 185350
rect 244942 185262 245122 185350
rect 245230 185262 245410 185350
rect 245664 185262 245844 185350
rect 245952 185262 246132 185350
rect 246240 185262 246420 185350
rect 246528 185262 246708 185350
rect 246816 185262 246996 185350
rect 247104 185262 247284 185350
rect 247392 185262 247572 185350
rect 247680 185262 247860 185350
rect 248114 185262 248294 185350
rect 248402 185262 248582 185350
rect 248690 185262 248870 185350
rect 248978 185262 249158 185350
rect 249266 185262 249446 185350
rect 249554 185262 249734 185350
rect 249842 185262 250022 185350
rect 250130 185262 250310 185350
rect 250564 185262 250744 185350
rect 360436 185262 360560 185350
rect 360814 185262 360994 185350
rect 361102 185262 361282 185350
rect 361390 185262 361570 185350
rect 361678 185262 361858 185350
rect 361966 185262 362146 185350
rect 362254 185262 362434 185350
rect 362542 185262 362722 185350
rect 362830 185262 363010 185350
rect 363264 185262 363444 185350
rect 363552 185262 363732 185350
rect 363840 185262 364020 185350
rect 364128 185262 364308 185350
rect 364416 185262 364596 185350
rect 364704 185262 364884 185350
rect 364992 185262 365172 185350
rect 365280 185262 365460 185350
rect 365714 185262 365894 185350
rect 366002 185262 366182 185350
rect 366290 185262 366470 185350
rect 366578 185262 366758 185350
rect 366866 185262 367046 185350
rect 367154 185262 367334 185350
rect 367442 185262 367622 185350
rect 367730 185262 367910 185350
rect 243214 184788 243394 184876
rect 243502 184788 243682 184876
rect 243790 184788 243970 184876
rect 244078 184788 244258 184876
rect 244366 184788 244546 184876
rect 244654 184788 244834 184876
rect 244942 184788 245122 184876
rect 245230 184788 245410 184876
rect 245664 184788 245844 184876
rect 245952 184788 246132 184876
rect 246240 184788 246420 184876
rect 246528 184788 246708 184876
rect 246816 184788 246996 184876
rect 247104 184788 247284 184876
rect 247392 184788 247572 184876
rect 247680 184788 247860 184876
rect 248114 184788 248294 184876
rect 248402 184788 248582 184876
rect 248690 184788 248870 184876
rect 248978 184788 249158 184876
rect 249266 184788 249446 184876
rect 249554 184788 249734 184876
rect 249842 184788 250022 184876
rect 250130 184788 250310 184876
rect 250564 184788 250744 184876
rect 360436 184788 360560 184876
rect 360814 184788 360994 184876
rect 361102 184788 361282 184876
rect 361390 184788 361570 184876
rect 361678 184788 361858 184876
rect 361966 184788 362146 184876
rect 362254 184788 362434 184876
rect 362542 184788 362722 184876
rect 362830 184788 363010 184876
rect 363264 184788 363444 184876
rect 363552 184788 363732 184876
rect 363840 184788 364020 184876
rect 364128 184788 364308 184876
rect 364416 184788 364596 184876
rect 364704 184788 364884 184876
rect 364992 184788 365172 184876
rect 365280 184788 365460 184876
rect 365714 184788 365894 184876
rect 366002 184788 366182 184876
rect 366290 184788 366470 184876
rect 366578 184788 366758 184876
rect 366866 184788 367046 184876
rect 367154 184788 367334 184876
rect 367442 184788 367622 184876
rect 367730 184788 367910 184876
rect 243214 184312 243394 184400
rect 243502 184312 243682 184400
rect 243790 184312 243970 184400
rect 244078 184312 244258 184400
rect 244366 184312 244546 184400
rect 244654 184312 244834 184400
rect 244942 184312 245122 184400
rect 245230 184312 245410 184400
rect 245664 184312 245844 184400
rect 245952 184312 246132 184400
rect 246240 184312 246420 184400
rect 246528 184312 246708 184400
rect 246816 184312 246996 184400
rect 247104 184312 247284 184400
rect 247392 184312 247572 184400
rect 247680 184312 247860 184400
rect 248114 184312 248294 184400
rect 248402 184312 248582 184400
rect 248690 184312 248870 184400
rect 248978 184312 249158 184400
rect 249266 184312 249446 184400
rect 249554 184312 249734 184400
rect 249842 184312 250022 184400
rect 250130 184312 250310 184400
rect 250564 184312 250744 184400
rect 360436 184312 360560 184400
rect 360814 184312 360994 184400
rect 361102 184312 361282 184400
rect 361390 184312 361570 184400
rect 361678 184312 361858 184400
rect 361966 184312 362146 184400
rect 362254 184312 362434 184400
rect 362542 184312 362722 184400
rect 362830 184312 363010 184400
rect 363264 184312 363444 184400
rect 363552 184312 363732 184400
rect 363840 184312 364020 184400
rect 364128 184312 364308 184400
rect 364416 184312 364596 184400
rect 364704 184312 364884 184400
rect 364992 184312 365172 184400
rect 365280 184312 365460 184400
rect 365714 184312 365894 184400
rect 366002 184312 366182 184400
rect 366290 184312 366470 184400
rect 366578 184312 366758 184400
rect 366866 184312 367046 184400
rect 367154 184312 367334 184400
rect 367442 184312 367622 184400
rect 367730 184312 367910 184400
rect 243214 184096 243394 184184
rect 243502 184096 243682 184184
rect 243790 184096 243970 184184
rect 244078 184096 244258 184184
rect 244366 184096 244546 184184
rect 244654 184096 244834 184184
rect 244942 184096 245122 184184
rect 245230 184096 245410 184184
rect 245664 184096 245844 184184
rect 245952 184096 246132 184184
rect 246240 184096 246420 184184
rect 246528 184096 246708 184184
rect 246816 184096 246996 184184
rect 247104 184096 247284 184184
rect 247392 184096 247572 184184
rect 247680 184096 247860 184184
rect 248114 184096 248294 184184
rect 248402 184096 248582 184184
rect 248690 184096 248870 184184
rect 248978 184096 249158 184184
rect 249266 184096 249446 184184
rect 249554 184096 249734 184184
rect 249842 184096 250022 184184
rect 250130 184096 250310 184184
rect 250564 184096 250744 184184
rect 360436 184096 360560 184184
rect 360814 184096 360994 184184
rect 361102 184096 361282 184184
rect 361390 184096 361570 184184
rect 361678 184096 361858 184184
rect 361966 184096 362146 184184
rect 362254 184096 362434 184184
rect 362542 184096 362722 184184
rect 362830 184096 363010 184184
rect 363264 184096 363444 184184
rect 363552 184096 363732 184184
rect 363840 184096 364020 184184
rect 364128 184096 364308 184184
rect 364416 184096 364596 184184
rect 364704 184096 364884 184184
rect 364992 184096 365172 184184
rect 365280 184096 365460 184184
rect 365714 184096 365894 184184
rect 366002 184096 366182 184184
rect 366290 184096 366470 184184
rect 366578 184096 366758 184184
rect 366866 184096 367046 184184
rect 367154 184096 367334 184184
rect 367442 184096 367622 184184
rect 367730 184096 367910 184184
rect 243214 183620 243394 183708
rect 243502 183620 243682 183708
rect 243790 183620 243970 183708
rect 244078 183620 244258 183708
rect 244366 183620 244546 183708
rect 244654 183620 244834 183708
rect 244942 183620 245122 183708
rect 245230 183620 245410 183708
rect 245664 183620 245844 183708
rect 245952 183620 246132 183708
rect 246240 183620 246420 183708
rect 246528 183620 246708 183708
rect 246816 183620 246996 183708
rect 247104 183620 247284 183708
rect 247392 183620 247572 183708
rect 247680 183620 247860 183708
rect 248114 183620 248294 183708
rect 248402 183620 248582 183708
rect 248690 183620 248870 183708
rect 248978 183620 249158 183708
rect 249266 183620 249446 183708
rect 249554 183620 249734 183708
rect 249842 183620 250022 183708
rect 250130 183620 250310 183708
rect 250564 183620 250744 183708
rect 360436 183620 360560 183708
rect 360814 183620 360994 183708
rect 361102 183620 361282 183708
rect 361390 183620 361570 183708
rect 361678 183620 361858 183708
rect 361966 183620 362146 183708
rect 362254 183620 362434 183708
rect 362542 183620 362722 183708
rect 362830 183620 363010 183708
rect 363264 183620 363444 183708
rect 363552 183620 363732 183708
rect 363840 183620 364020 183708
rect 364128 183620 364308 183708
rect 364416 183620 364596 183708
rect 364704 183620 364884 183708
rect 364992 183620 365172 183708
rect 365280 183620 365460 183708
rect 365714 183620 365894 183708
rect 366002 183620 366182 183708
rect 366290 183620 366470 183708
rect 366578 183620 366758 183708
rect 366866 183620 367046 183708
rect 367154 183620 367334 183708
rect 367442 183620 367622 183708
rect 367730 183620 367910 183708
rect 243214 183404 243394 183492
rect 243502 183404 243682 183492
rect 243790 183404 243970 183492
rect 244078 183404 244258 183492
rect 244366 183404 244546 183492
rect 244654 183404 244834 183492
rect 244942 183404 245122 183492
rect 245230 183404 245410 183492
rect 245664 183404 245844 183492
rect 245952 183404 246132 183492
rect 246240 183404 246420 183492
rect 246528 183404 246708 183492
rect 246816 183404 246996 183492
rect 247104 183404 247284 183492
rect 247392 183404 247572 183492
rect 247680 183404 247860 183492
rect 248114 183404 248294 183492
rect 248402 183404 248582 183492
rect 248690 183404 248870 183492
rect 248978 183404 249158 183492
rect 249266 183404 249446 183492
rect 249554 183404 249734 183492
rect 249842 183404 250022 183492
rect 250130 183404 250310 183492
rect 250564 183404 250744 183492
rect 360436 183404 360560 183492
rect 360814 183404 360994 183492
rect 361102 183404 361282 183492
rect 361390 183404 361570 183492
rect 361678 183404 361858 183492
rect 361966 183404 362146 183492
rect 362254 183404 362434 183492
rect 362542 183404 362722 183492
rect 362830 183404 363010 183492
rect 363264 183404 363444 183492
rect 363552 183404 363732 183492
rect 363840 183404 364020 183492
rect 364128 183404 364308 183492
rect 364416 183404 364596 183492
rect 364704 183404 364884 183492
rect 364992 183404 365172 183492
rect 365280 183404 365460 183492
rect 365714 183404 365894 183492
rect 366002 183404 366182 183492
rect 366290 183404 366470 183492
rect 366578 183404 366758 183492
rect 366866 183404 367046 183492
rect 367154 183404 367334 183492
rect 367442 183404 367622 183492
rect 367730 183404 367910 183492
rect 243214 182928 243394 183016
rect 243502 182928 243682 183016
rect 243790 182928 243970 183016
rect 244078 182928 244258 183016
rect 244366 182928 244546 183016
rect 244654 182928 244834 183016
rect 244942 182928 245122 183016
rect 245230 182928 245410 183016
rect 245664 182928 245844 183016
rect 245952 182928 246132 183016
rect 246240 182928 246420 183016
rect 246528 182928 246708 183016
rect 246816 182928 246996 183016
rect 247104 182928 247284 183016
rect 247392 182928 247572 183016
rect 247680 182928 247860 183016
rect 248114 182928 248294 183016
rect 248402 182928 248582 183016
rect 248690 182928 248870 183016
rect 248978 182928 249158 183016
rect 249266 182928 249446 183016
rect 249554 182928 249734 183016
rect 249842 182928 250022 183016
rect 250130 182928 250310 183016
rect 250564 182928 250744 183016
rect 360436 182928 360560 183016
rect 360814 182928 360994 183016
rect 361102 182928 361282 183016
rect 361390 182928 361570 183016
rect 361678 182928 361858 183016
rect 361966 182928 362146 183016
rect 362254 182928 362434 183016
rect 362542 182928 362722 183016
rect 362830 182928 363010 183016
rect 363264 182928 363444 183016
rect 363552 182928 363732 183016
rect 363840 182928 364020 183016
rect 364128 182928 364308 183016
rect 364416 182928 364596 183016
rect 364704 182928 364884 183016
rect 364992 182928 365172 183016
rect 365280 182928 365460 183016
rect 365714 182928 365894 183016
rect 366002 182928 366182 183016
rect 366290 182928 366470 183016
rect 366578 182928 366758 183016
rect 366866 182928 367046 183016
rect 367154 182928 367334 183016
rect 367442 182928 367622 183016
rect 367730 182928 367910 183016
rect 243214 182712 243394 182800
rect 243502 182712 243682 182800
rect 243790 182712 243970 182800
rect 244078 182712 244258 182800
rect 244366 182712 244546 182800
rect 244654 182712 244834 182800
rect 244942 182712 245122 182800
rect 245230 182712 245410 182800
rect 245664 182712 245844 182800
rect 245952 182712 246132 182800
rect 246240 182712 246420 182800
rect 246528 182712 246708 182800
rect 246816 182712 246996 182800
rect 247104 182712 247284 182800
rect 247392 182712 247572 182800
rect 247680 182712 247860 182800
rect 248114 182712 248294 182800
rect 248402 182712 248582 182800
rect 248690 182712 248870 182800
rect 248978 182712 249158 182800
rect 249266 182712 249446 182800
rect 249554 182712 249734 182800
rect 249842 182712 250022 182800
rect 250130 182712 250310 182800
rect 250564 182712 250744 182800
rect 360436 182712 360560 182800
rect 360814 182712 360994 182800
rect 361102 182712 361282 182800
rect 361390 182712 361570 182800
rect 361678 182712 361858 182800
rect 361966 182712 362146 182800
rect 362254 182712 362434 182800
rect 362542 182712 362722 182800
rect 362830 182712 363010 182800
rect 363264 182712 363444 182800
rect 363552 182712 363732 182800
rect 363840 182712 364020 182800
rect 364128 182712 364308 182800
rect 364416 182712 364596 182800
rect 364704 182712 364884 182800
rect 364992 182712 365172 182800
rect 365280 182712 365460 182800
rect 365714 182712 365894 182800
rect 366002 182712 366182 182800
rect 366290 182712 366470 182800
rect 366578 182712 366758 182800
rect 366866 182712 367046 182800
rect 367154 182712 367334 182800
rect 367442 182712 367622 182800
rect 367730 182712 367910 182800
rect 243214 182236 243394 182324
rect 243502 182236 243682 182324
rect 243790 182236 243970 182324
rect 244078 182236 244258 182324
rect 244366 182236 244546 182324
rect 244654 182236 244834 182324
rect 244942 182236 245122 182324
rect 245230 182236 245410 182324
rect 245664 182236 245844 182324
rect 245952 182236 246132 182324
rect 246240 182236 246420 182324
rect 246528 182236 246708 182324
rect 246816 182236 246996 182324
rect 247104 182236 247284 182324
rect 247392 182236 247572 182324
rect 247680 182236 247860 182324
rect 248114 182236 248294 182324
rect 248402 182236 248582 182324
rect 248690 182236 248870 182324
rect 248978 182236 249158 182324
rect 249266 182236 249446 182324
rect 249554 182236 249734 182324
rect 249842 182236 250022 182324
rect 250130 182236 250310 182324
rect 250564 182236 250744 182324
rect 360436 182236 360560 182324
rect 360814 182236 360994 182324
rect 361102 182236 361282 182324
rect 361390 182236 361570 182324
rect 361678 182236 361858 182324
rect 361966 182236 362146 182324
rect 362254 182236 362434 182324
rect 362542 182236 362722 182324
rect 362830 182236 363010 182324
rect 363264 182236 363444 182324
rect 363552 182236 363732 182324
rect 363840 182236 364020 182324
rect 364128 182236 364308 182324
rect 364416 182236 364596 182324
rect 364704 182236 364884 182324
rect 364992 182236 365172 182324
rect 365280 182236 365460 182324
rect 365714 182236 365894 182324
rect 366002 182236 366182 182324
rect 366290 182236 366470 182324
rect 366578 182236 366758 182324
rect 366866 182236 367046 182324
rect 367154 182236 367334 182324
rect 367442 182236 367622 182324
rect 367730 182236 367910 182324
rect 243214 181762 243394 181850
rect 243502 181762 243682 181850
rect 243790 181762 243970 181850
rect 244078 181762 244258 181850
rect 244366 181762 244546 181850
rect 244654 181762 244834 181850
rect 244942 181762 245122 181850
rect 245230 181762 245410 181850
rect 245664 181762 245844 181850
rect 245952 181762 246132 181850
rect 246240 181762 246420 181850
rect 246528 181762 246708 181850
rect 246816 181762 246996 181850
rect 247104 181762 247284 181850
rect 247392 181762 247572 181850
rect 247680 181762 247860 181850
rect 248114 181762 248294 181850
rect 248402 181762 248582 181850
rect 248690 181762 248870 181850
rect 248978 181762 249158 181850
rect 249266 181762 249446 181850
rect 249554 181762 249734 181850
rect 249842 181762 250022 181850
rect 250130 181762 250310 181850
rect 250564 181762 250744 181850
rect 360436 181762 360560 181850
rect 360814 181762 360994 181850
rect 361102 181762 361282 181850
rect 361390 181762 361570 181850
rect 361678 181762 361858 181850
rect 361966 181762 362146 181850
rect 362254 181762 362434 181850
rect 362542 181762 362722 181850
rect 362830 181762 363010 181850
rect 363264 181762 363444 181850
rect 363552 181762 363732 181850
rect 363840 181762 364020 181850
rect 364128 181762 364308 181850
rect 364416 181762 364596 181850
rect 364704 181762 364884 181850
rect 364992 181762 365172 181850
rect 365280 181762 365460 181850
rect 365714 181762 365894 181850
rect 366002 181762 366182 181850
rect 366290 181762 366470 181850
rect 366578 181762 366758 181850
rect 366866 181762 367046 181850
rect 367154 181762 367334 181850
rect 367442 181762 367622 181850
rect 367730 181762 367910 181850
rect 243214 181286 243394 181374
rect 243502 181286 243682 181374
rect 243790 181286 243970 181374
rect 244078 181286 244258 181374
rect 244366 181286 244546 181374
rect 244654 181286 244834 181374
rect 244942 181286 245122 181374
rect 245230 181286 245410 181374
rect 245664 181286 245844 181374
rect 245952 181286 246132 181374
rect 246240 181286 246420 181374
rect 246528 181286 246708 181374
rect 246816 181286 246996 181374
rect 247104 181286 247284 181374
rect 247392 181286 247572 181374
rect 247680 181286 247860 181374
rect 248114 181286 248294 181374
rect 248402 181286 248582 181374
rect 248690 181286 248870 181374
rect 248978 181286 249158 181374
rect 249266 181286 249446 181374
rect 249554 181286 249734 181374
rect 249842 181286 250022 181374
rect 250130 181286 250310 181374
rect 250564 181286 250744 181374
rect 360436 181286 360560 181374
rect 360814 181286 360994 181374
rect 361102 181286 361282 181374
rect 361390 181286 361570 181374
rect 361678 181286 361858 181374
rect 361966 181286 362146 181374
rect 362254 181286 362434 181374
rect 362542 181286 362722 181374
rect 362830 181286 363010 181374
rect 363264 181286 363444 181374
rect 363552 181286 363732 181374
rect 363840 181286 364020 181374
rect 364128 181286 364308 181374
rect 364416 181286 364596 181374
rect 364704 181286 364884 181374
rect 364992 181286 365172 181374
rect 365280 181286 365460 181374
rect 365714 181286 365894 181374
rect 366002 181286 366182 181374
rect 366290 181286 366470 181374
rect 366578 181286 366758 181374
rect 366866 181286 367046 181374
rect 367154 181286 367334 181374
rect 367442 181286 367622 181374
rect 367730 181286 367910 181374
rect 243214 181070 243394 181158
rect 243502 181070 243682 181158
rect 243790 181070 243970 181158
rect 244078 181070 244258 181158
rect 244366 181070 244546 181158
rect 244654 181070 244834 181158
rect 244942 181070 245122 181158
rect 245230 181070 245410 181158
rect 245664 181070 245844 181158
rect 245952 181070 246132 181158
rect 246240 181070 246420 181158
rect 246528 181070 246708 181158
rect 246816 181070 246996 181158
rect 247104 181070 247284 181158
rect 247392 181070 247572 181158
rect 247680 181070 247860 181158
rect 248114 181070 248294 181158
rect 248402 181070 248582 181158
rect 248690 181070 248870 181158
rect 248978 181070 249158 181158
rect 249266 181070 249446 181158
rect 249554 181070 249734 181158
rect 249842 181070 250022 181158
rect 250130 181070 250310 181158
rect 250564 181070 250744 181158
rect 360436 181070 360560 181158
rect 360814 181070 360994 181158
rect 361102 181070 361282 181158
rect 361390 181070 361570 181158
rect 361678 181070 361858 181158
rect 361966 181070 362146 181158
rect 362254 181070 362434 181158
rect 362542 181070 362722 181158
rect 362830 181070 363010 181158
rect 363264 181070 363444 181158
rect 363552 181070 363732 181158
rect 363840 181070 364020 181158
rect 364128 181070 364308 181158
rect 364416 181070 364596 181158
rect 364704 181070 364884 181158
rect 364992 181070 365172 181158
rect 365280 181070 365460 181158
rect 365714 181070 365894 181158
rect 366002 181070 366182 181158
rect 366290 181070 366470 181158
rect 366578 181070 366758 181158
rect 366866 181070 367046 181158
rect 367154 181070 367334 181158
rect 367442 181070 367622 181158
rect 367730 181070 367910 181158
rect 243214 180594 243394 180682
rect 243502 180594 243682 180682
rect 243790 180594 243970 180682
rect 244078 180594 244258 180682
rect 244366 180594 244546 180682
rect 244654 180594 244834 180682
rect 244942 180594 245122 180682
rect 245230 180594 245410 180682
rect 245664 180594 245844 180682
rect 245952 180594 246132 180682
rect 246240 180594 246420 180682
rect 246528 180594 246708 180682
rect 246816 180594 246996 180682
rect 247104 180594 247284 180682
rect 247392 180594 247572 180682
rect 247680 180594 247860 180682
rect 248114 180594 248294 180682
rect 248402 180594 248582 180682
rect 248690 180594 248870 180682
rect 248978 180594 249158 180682
rect 249266 180594 249446 180682
rect 249554 180594 249734 180682
rect 249842 180594 250022 180682
rect 250130 180594 250310 180682
rect 250564 180594 250744 180682
rect 360436 180594 360560 180682
rect 360814 180594 360994 180682
rect 361102 180594 361282 180682
rect 361390 180594 361570 180682
rect 361678 180594 361858 180682
rect 361966 180594 362146 180682
rect 362254 180594 362434 180682
rect 362542 180594 362722 180682
rect 362830 180594 363010 180682
rect 363264 180594 363444 180682
rect 363552 180594 363732 180682
rect 363840 180594 364020 180682
rect 364128 180594 364308 180682
rect 364416 180594 364596 180682
rect 364704 180594 364884 180682
rect 364992 180594 365172 180682
rect 365280 180594 365460 180682
rect 365714 180594 365894 180682
rect 366002 180594 366182 180682
rect 366290 180594 366470 180682
rect 366578 180594 366758 180682
rect 366866 180594 367046 180682
rect 367154 180594 367334 180682
rect 367442 180594 367622 180682
rect 367730 180594 367910 180682
rect 243214 180378 243394 180466
rect 243502 180378 243682 180466
rect 243790 180378 243970 180466
rect 244078 180378 244258 180466
rect 244366 180378 244546 180466
rect 244654 180378 244834 180466
rect 244942 180378 245122 180466
rect 245230 180378 245410 180466
rect 245664 180378 245844 180466
rect 245952 180378 246132 180466
rect 246240 180378 246420 180466
rect 246528 180378 246708 180466
rect 246816 180378 246996 180466
rect 247104 180378 247284 180466
rect 247392 180378 247572 180466
rect 247680 180378 247860 180466
rect 248114 180378 248294 180466
rect 248402 180378 248582 180466
rect 248690 180378 248870 180466
rect 248978 180378 249158 180466
rect 249266 180378 249446 180466
rect 249554 180378 249734 180466
rect 249842 180378 250022 180466
rect 250130 180378 250310 180466
rect 250564 180378 250744 180466
rect 360436 180378 360560 180466
rect 360814 180378 360994 180466
rect 361102 180378 361282 180466
rect 361390 180378 361570 180466
rect 361678 180378 361858 180466
rect 361966 180378 362146 180466
rect 362254 180378 362434 180466
rect 362542 180378 362722 180466
rect 362830 180378 363010 180466
rect 363264 180378 363444 180466
rect 363552 180378 363732 180466
rect 363840 180378 364020 180466
rect 364128 180378 364308 180466
rect 364416 180378 364596 180466
rect 364704 180378 364884 180466
rect 364992 180378 365172 180466
rect 365280 180378 365460 180466
rect 365714 180378 365894 180466
rect 366002 180378 366182 180466
rect 366290 180378 366470 180466
rect 366578 180378 366758 180466
rect 366866 180378 367046 180466
rect 367154 180378 367334 180466
rect 367442 180378 367622 180466
rect 367730 180378 367910 180466
rect 243214 179902 243394 179990
rect 243502 179902 243682 179990
rect 243790 179902 243970 179990
rect 244078 179902 244258 179990
rect 244366 179902 244546 179990
rect 244654 179902 244834 179990
rect 244942 179902 245122 179990
rect 245230 179902 245410 179990
rect 245664 179902 245844 179990
rect 245952 179902 246132 179990
rect 246240 179902 246420 179990
rect 246528 179902 246708 179990
rect 246816 179902 246996 179990
rect 247104 179902 247284 179990
rect 247392 179902 247572 179990
rect 247680 179902 247860 179990
rect 248114 179902 248294 179990
rect 248402 179902 248582 179990
rect 248690 179902 248870 179990
rect 248978 179902 249158 179990
rect 249266 179902 249446 179990
rect 249554 179902 249734 179990
rect 249842 179902 250022 179990
rect 250130 179902 250310 179990
rect 250564 179902 250744 179990
rect 360436 179902 360560 179990
rect 360814 179902 360994 179990
rect 361102 179902 361282 179990
rect 361390 179902 361570 179990
rect 361678 179902 361858 179990
rect 361966 179902 362146 179990
rect 362254 179902 362434 179990
rect 362542 179902 362722 179990
rect 362830 179902 363010 179990
rect 363264 179902 363444 179990
rect 363552 179902 363732 179990
rect 363840 179902 364020 179990
rect 364128 179902 364308 179990
rect 364416 179902 364596 179990
rect 364704 179902 364884 179990
rect 364992 179902 365172 179990
rect 365280 179902 365460 179990
rect 365714 179902 365894 179990
rect 366002 179902 366182 179990
rect 366290 179902 366470 179990
rect 366578 179902 366758 179990
rect 366866 179902 367046 179990
rect 367154 179902 367334 179990
rect 367442 179902 367622 179990
rect 367730 179902 367910 179990
rect 243214 179686 243394 179774
rect 243502 179686 243682 179774
rect 243790 179686 243970 179774
rect 244078 179686 244258 179774
rect 244366 179686 244546 179774
rect 244654 179686 244834 179774
rect 244942 179686 245122 179774
rect 245230 179686 245410 179774
rect 245664 179686 245844 179774
rect 245952 179686 246132 179774
rect 246240 179686 246420 179774
rect 246528 179686 246708 179774
rect 246816 179686 246996 179774
rect 247104 179686 247284 179774
rect 247392 179686 247572 179774
rect 247680 179686 247860 179774
rect 248114 179686 248294 179774
rect 248402 179686 248582 179774
rect 248690 179686 248870 179774
rect 248978 179686 249158 179774
rect 249266 179686 249446 179774
rect 249554 179686 249734 179774
rect 249842 179686 250022 179774
rect 250130 179686 250310 179774
rect 250564 179686 250744 179774
rect 360436 179686 360560 179774
rect 360814 179686 360994 179774
rect 361102 179686 361282 179774
rect 361390 179686 361570 179774
rect 361678 179686 361858 179774
rect 361966 179686 362146 179774
rect 362254 179686 362434 179774
rect 362542 179686 362722 179774
rect 362830 179686 363010 179774
rect 363264 179686 363444 179774
rect 363552 179686 363732 179774
rect 363840 179686 364020 179774
rect 364128 179686 364308 179774
rect 364416 179686 364596 179774
rect 364704 179686 364884 179774
rect 364992 179686 365172 179774
rect 365280 179686 365460 179774
rect 365714 179686 365894 179774
rect 366002 179686 366182 179774
rect 366290 179686 366470 179774
rect 366578 179686 366758 179774
rect 366866 179686 367046 179774
rect 367154 179686 367334 179774
rect 367442 179686 367622 179774
rect 367730 179686 367910 179774
rect 243214 179210 243394 179298
rect 243502 179210 243682 179298
rect 243790 179210 243970 179298
rect 244078 179210 244258 179298
rect 244366 179210 244546 179298
rect 244654 179210 244834 179298
rect 244942 179210 245122 179298
rect 245230 179210 245410 179298
rect 245664 179210 245844 179298
rect 245952 179210 246132 179298
rect 246240 179210 246420 179298
rect 246528 179210 246708 179298
rect 246816 179210 246996 179298
rect 247104 179210 247284 179298
rect 247392 179210 247572 179298
rect 247680 179210 247860 179298
rect 248114 179210 248294 179298
rect 248402 179210 248582 179298
rect 248690 179210 248870 179298
rect 248978 179210 249158 179298
rect 249266 179210 249446 179298
rect 249554 179210 249734 179298
rect 249842 179210 250022 179298
rect 250130 179210 250310 179298
rect 250564 179210 250744 179298
rect 360436 179210 360560 179298
rect 360814 179210 360994 179298
rect 361102 179210 361282 179298
rect 361390 179210 361570 179298
rect 361678 179210 361858 179298
rect 361966 179210 362146 179298
rect 362254 179210 362434 179298
rect 362542 179210 362722 179298
rect 362830 179210 363010 179298
rect 363264 179210 363444 179298
rect 363552 179210 363732 179298
rect 363840 179210 364020 179298
rect 364128 179210 364308 179298
rect 364416 179210 364596 179298
rect 364704 179210 364884 179298
rect 364992 179210 365172 179298
rect 365280 179210 365460 179298
rect 365714 179210 365894 179298
rect 366002 179210 366182 179298
rect 366290 179210 366470 179298
rect 366578 179210 366758 179298
rect 366866 179210 367046 179298
rect 367154 179210 367334 179298
rect 367442 179210 367622 179298
rect 367730 179210 367910 179298
rect 243214 178736 243394 178824
rect 243502 178736 243682 178824
rect 243790 178736 243970 178824
rect 244078 178736 244258 178824
rect 244366 178736 244546 178824
rect 244654 178736 244834 178824
rect 244942 178736 245122 178824
rect 245230 178736 245410 178824
rect 245664 178736 245844 178824
rect 245952 178736 246132 178824
rect 246240 178736 246420 178824
rect 246528 178736 246708 178824
rect 246816 178736 246996 178824
rect 247104 178736 247284 178824
rect 247392 178736 247572 178824
rect 247680 178736 247860 178824
rect 248114 178736 248294 178824
rect 248402 178736 248582 178824
rect 248690 178736 248870 178824
rect 248978 178736 249158 178824
rect 249266 178736 249446 178824
rect 249554 178736 249734 178824
rect 249842 178736 250022 178824
rect 250130 178736 250310 178824
rect 250564 178736 250744 178824
rect 360436 178736 360560 178824
rect 360814 178736 360994 178824
rect 361102 178736 361282 178824
rect 361390 178736 361570 178824
rect 361678 178736 361858 178824
rect 361966 178736 362146 178824
rect 362254 178736 362434 178824
rect 362542 178736 362722 178824
rect 362830 178736 363010 178824
rect 363264 178736 363444 178824
rect 363552 178736 363732 178824
rect 363840 178736 364020 178824
rect 364128 178736 364308 178824
rect 364416 178736 364596 178824
rect 364704 178736 364884 178824
rect 364992 178736 365172 178824
rect 365280 178736 365460 178824
rect 365714 178736 365894 178824
rect 366002 178736 366182 178824
rect 366290 178736 366470 178824
rect 366578 178736 366758 178824
rect 366866 178736 367046 178824
rect 367154 178736 367334 178824
rect 367442 178736 367622 178824
rect 367730 178736 367910 178824
rect 243214 178260 243394 178348
rect 243502 178260 243682 178348
rect 243790 178260 243970 178348
rect 244078 178260 244258 178348
rect 244366 178260 244546 178348
rect 244654 178260 244834 178348
rect 244942 178260 245122 178348
rect 245230 178260 245410 178348
rect 245664 178260 245844 178348
rect 245952 178260 246132 178348
rect 246240 178260 246420 178348
rect 246528 178260 246708 178348
rect 246816 178260 246996 178348
rect 247104 178260 247284 178348
rect 247392 178260 247572 178348
rect 247680 178260 247860 178348
rect 248114 178260 248294 178348
rect 248402 178260 248582 178348
rect 248690 178260 248870 178348
rect 248978 178260 249158 178348
rect 249266 178260 249446 178348
rect 249554 178260 249734 178348
rect 249842 178260 250022 178348
rect 250130 178260 250310 178348
rect 250564 178260 250744 178348
rect 360436 178260 360560 178348
rect 360814 178260 360994 178348
rect 361102 178260 361282 178348
rect 361390 178260 361570 178348
rect 361678 178260 361858 178348
rect 361966 178260 362146 178348
rect 362254 178260 362434 178348
rect 362542 178260 362722 178348
rect 362830 178260 363010 178348
rect 363264 178260 363444 178348
rect 363552 178260 363732 178348
rect 363840 178260 364020 178348
rect 364128 178260 364308 178348
rect 364416 178260 364596 178348
rect 364704 178260 364884 178348
rect 364992 178260 365172 178348
rect 365280 178260 365460 178348
rect 365714 178260 365894 178348
rect 366002 178260 366182 178348
rect 366290 178260 366470 178348
rect 366578 178260 366758 178348
rect 366866 178260 367046 178348
rect 367154 178260 367334 178348
rect 367442 178260 367622 178348
rect 367730 178260 367910 178348
rect 243214 178044 243394 178132
rect 243502 178044 243682 178132
rect 243790 178044 243970 178132
rect 244078 178044 244258 178132
rect 244366 178044 244546 178132
rect 244654 178044 244834 178132
rect 244942 178044 245122 178132
rect 245230 178044 245410 178132
rect 245664 178044 245844 178132
rect 245952 178044 246132 178132
rect 246240 178044 246420 178132
rect 246528 178044 246708 178132
rect 246816 178044 246996 178132
rect 247104 178044 247284 178132
rect 247392 178044 247572 178132
rect 247680 178044 247860 178132
rect 248114 178044 248294 178132
rect 248402 178044 248582 178132
rect 248690 178044 248870 178132
rect 248978 178044 249158 178132
rect 249266 178044 249446 178132
rect 249554 178044 249734 178132
rect 249842 178044 250022 178132
rect 250130 178044 250310 178132
rect 250564 178044 250744 178132
rect 360436 178044 360560 178132
rect 360814 178044 360994 178132
rect 361102 178044 361282 178132
rect 361390 178044 361570 178132
rect 361678 178044 361858 178132
rect 361966 178044 362146 178132
rect 362254 178044 362434 178132
rect 362542 178044 362722 178132
rect 362830 178044 363010 178132
rect 363264 178044 363444 178132
rect 363552 178044 363732 178132
rect 363840 178044 364020 178132
rect 364128 178044 364308 178132
rect 364416 178044 364596 178132
rect 364704 178044 364884 178132
rect 364992 178044 365172 178132
rect 365280 178044 365460 178132
rect 365714 178044 365894 178132
rect 366002 178044 366182 178132
rect 366290 178044 366470 178132
rect 366578 178044 366758 178132
rect 366866 178044 367046 178132
rect 367154 178044 367334 178132
rect 367442 178044 367622 178132
rect 367730 178044 367910 178132
rect 243214 177568 243394 177656
rect 243502 177568 243682 177656
rect 243790 177568 243970 177656
rect 244078 177568 244258 177656
rect 244366 177568 244546 177656
rect 244654 177568 244834 177656
rect 244942 177568 245122 177656
rect 245230 177568 245410 177656
rect 245664 177568 245844 177656
rect 245952 177568 246132 177656
rect 246240 177568 246420 177656
rect 246528 177568 246708 177656
rect 246816 177568 246996 177656
rect 247104 177568 247284 177656
rect 247392 177568 247572 177656
rect 247680 177568 247860 177656
rect 248114 177568 248294 177656
rect 248402 177568 248582 177656
rect 248690 177568 248870 177656
rect 248978 177568 249158 177656
rect 249266 177568 249446 177656
rect 249554 177568 249734 177656
rect 249842 177568 250022 177656
rect 250130 177568 250310 177656
rect 250564 177568 250744 177656
rect 360436 177568 360560 177656
rect 360814 177568 360994 177656
rect 361102 177568 361282 177656
rect 361390 177568 361570 177656
rect 361678 177568 361858 177656
rect 361966 177568 362146 177656
rect 362254 177568 362434 177656
rect 362542 177568 362722 177656
rect 362830 177568 363010 177656
rect 363264 177568 363444 177656
rect 363552 177568 363732 177656
rect 363840 177568 364020 177656
rect 364128 177568 364308 177656
rect 364416 177568 364596 177656
rect 364704 177568 364884 177656
rect 364992 177568 365172 177656
rect 365280 177568 365460 177656
rect 365714 177568 365894 177656
rect 366002 177568 366182 177656
rect 366290 177568 366470 177656
rect 366578 177568 366758 177656
rect 366866 177568 367046 177656
rect 367154 177568 367334 177656
rect 367442 177568 367622 177656
rect 367730 177568 367910 177656
rect 243214 177352 243394 177440
rect 243502 177352 243682 177440
rect 243790 177352 243970 177440
rect 244078 177352 244258 177440
rect 244366 177352 244546 177440
rect 244654 177352 244834 177440
rect 244942 177352 245122 177440
rect 245230 177352 245410 177440
rect 245664 177352 245844 177440
rect 245952 177352 246132 177440
rect 246240 177352 246420 177440
rect 246528 177352 246708 177440
rect 246816 177352 246996 177440
rect 247104 177352 247284 177440
rect 247392 177352 247572 177440
rect 247680 177352 247860 177440
rect 248114 177352 248294 177440
rect 248402 177352 248582 177440
rect 248690 177352 248870 177440
rect 248978 177352 249158 177440
rect 249266 177352 249446 177440
rect 249554 177352 249734 177440
rect 249842 177352 250022 177440
rect 250130 177352 250310 177440
rect 250564 177352 250744 177440
rect 360436 177352 360560 177440
rect 360814 177352 360994 177440
rect 361102 177352 361282 177440
rect 361390 177352 361570 177440
rect 361678 177352 361858 177440
rect 361966 177352 362146 177440
rect 362254 177352 362434 177440
rect 362542 177352 362722 177440
rect 362830 177352 363010 177440
rect 363264 177352 363444 177440
rect 363552 177352 363732 177440
rect 363840 177352 364020 177440
rect 364128 177352 364308 177440
rect 364416 177352 364596 177440
rect 364704 177352 364884 177440
rect 364992 177352 365172 177440
rect 365280 177352 365460 177440
rect 365714 177352 365894 177440
rect 366002 177352 366182 177440
rect 366290 177352 366470 177440
rect 366578 177352 366758 177440
rect 366866 177352 367046 177440
rect 367154 177352 367334 177440
rect 367442 177352 367622 177440
rect 367730 177352 367910 177440
rect 243214 176876 243394 176964
rect 243502 176876 243682 176964
rect 243790 176876 243970 176964
rect 244078 176876 244258 176964
rect 244366 176876 244546 176964
rect 244654 176876 244834 176964
rect 244942 176876 245122 176964
rect 245230 176876 245410 176964
rect 245664 176876 245844 176964
rect 245952 176876 246132 176964
rect 246240 176876 246420 176964
rect 246528 176876 246708 176964
rect 246816 176876 246996 176964
rect 247104 176876 247284 176964
rect 247392 176876 247572 176964
rect 247680 176876 247860 176964
rect 248114 176876 248294 176964
rect 248402 176876 248582 176964
rect 248690 176876 248870 176964
rect 248978 176876 249158 176964
rect 249266 176876 249446 176964
rect 249554 176876 249734 176964
rect 249842 176876 250022 176964
rect 250130 176876 250310 176964
rect 250564 176876 250744 176964
rect 360436 176876 360560 176964
rect 360814 176876 360994 176964
rect 361102 176876 361282 176964
rect 361390 176876 361570 176964
rect 361678 176876 361858 176964
rect 361966 176876 362146 176964
rect 362254 176876 362434 176964
rect 362542 176876 362722 176964
rect 362830 176876 363010 176964
rect 363264 176876 363444 176964
rect 363552 176876 363732 176964
rect 363840 176876 364020 176964
rect 364128 176876 364308 176964
rect 364416 176876 364596 176964
rect 364704 176876 364884 176964
rect 364992 176876 365172 176964
rect 365280 176876 365460 176964
rect 365714 176876 365894 176964
rect 366002 176876 366182 176964
rect 366290 176876 366470 176964
rect 366578 176876 366758 176964
rect 366866 176876 367046 176964
rect 367154 176876 367334 176964
rect 367442 176876 367622 176964
rect 367730 176876 367910 176964
rect 243214 176660 243394 176748
rect 243502 176660 243682 176748
rect 243790 176660 243970 176748
rect 244078 176660 244258 176748
rect 244366 176660 244546 176748
rect 244654 176660 244834 176748
rect 244942 176660 245122 176748
rect 245230 176660 245410 176748
rect 245664 176660 245844 176748
rect 245952 176660 246132 176748
rect 246240 176660 246420 176748
rect 246528 176660 246708 176748
rect 246816 176660 246996 176748
rect 247104 176660 247284 176748
rect 247392 176660 247572 176748
rect 247680 176660 247860 176748
rect 248114 176660 248294 176748
rect 248402 176660 248582 176748
rect 248690 176660 248870 176748
rect 248978 176660 249158 176748
rect 249266 176660 249446 176748
rect 249554 176660 249734 176748
rect 249842 176660 250022 176748
rect 250130 176660 250310 176748
rect 250564 176660 250744 176748
rect 360436 176660 360560 176748
rect 360814 176660 360994 176748
rect 361102 176660 361282 176748
rect 361390 176660 361570 176748
rect 361678 176660 361858 176748
rect 361966 176660 362146 176748
rect 362254 176660 362434 176748
rect 362542 176660 362722 176748
rect 362830 176660 363010 176748
rect 363264 176660 363444 176748
rect 363552 176660 363732 176748
rect 363840 176660 364020 176748
rect 364128 176660 364308 176748
rect 364416 176660 364596 176748
rect 364704 176660 364884 176748
rect 364992 176660 365172 176748
rect 365280 176660 365460 176748
rect 365714 176660 365894 176748
rect 366002 176660 366182 176748
rect 366290 176660 366470 176748
rect 366578 176660 366758 176748
rect 366866 176660 367046 176748
rect 367154 176660 367334 176748
rect 367442 176660 367622 176748
rect 367730 176660 367910 176748
rect 243214 176184 243394 176272
rect 243502 176184 243682 176272
rect 243790 176184 243970 176272
rect 244078 176184 244258 176272
rect 244366 176184 244546 176272
rect 244654 176184 244834 176272
rect 244942 176184 245122 176272
rect 245230 176184 245410 176272
rect 245664 176184 245844 176272
rect 245952 176184 246132 176272
rect 246240 176184 246420 176272
rect 246528 176184 246708 176272
rect 246816 176184 246996 176272
rect 247104 176184 247284 176272
rect 247392 176184 247572 176272
rect 247680 176184 247860 176272
rect 248114 176184 248294 176272
rect 248402 176184 248582 176272
rect 248690 176184 248870 176272
rect 248978 176184 249158 176272
rect 249266 176184 249446 176272
rect 249554 176184 249734 176272
rect 249842 176184 250022 176272
rect 250130 176184 250310 176272
rect 250564 176184 250744 176272
rect 360436 176184 360560 176272
rect 360814 176184 360994 176272
rect 361102 176184 361282 176272
rect 361390 176184 361570 176272
rect 361678 176184 361858 176272
rect 361966 176184 362146 176272
rect 362254 176184 362434 176272
rect 362542 176184 362722 176272
rect 362830 176184 363010 176272
rect 363264 176184 363444 176272
rect 363552 176184 363732 176272
rect 363840 176184 364020 176272
rect 364128 176184 364308 176272
rect 364416 176184 364596 176272
rect 364704 176184 364884 176272
rect 364992 176184 365172 176272
rect 365280 176184 365460 176272
rect 365714 176184 365894 176272
rect 366002 176184 366182 176272
rect 366290 176184 366470 176272
rect 366578 176184 366758 176272
rect 366866 176184 367046 176272
rect 367154 176184 367334 176272
rect 367442 176184 367622 176272
rect 367730 176184 367910 176272
rect 243214 175710 243394 175798
rect 243502 175710 243682 175798
rect 243790 175710 243970 175798
rect 244078 175710 244258 175798
rect 244366 175710 244546 175798
rect 244654 175710 244834 175798
rect 244942 175710 245122 175798
rect 245230 175710 245410 175798
rect 245664 175710 245844 175798
rect 245952 175710 246132 175798
rect 246240 175710 246420 175798
rect 246528 175710 246708 175798
rect 246816 175710 246996 175798
rect 247104 175710 247284 175798
rect 247392 175710 247572 175798
rect 247680 175710 247860 175798
rect 248114 175710 248294 175798
rect 248402 175710 248582 175798
rect 248690 175710 248870 175798
rect 248978 175710 249158 175798
rect 249266 175710 249446 175798
rect 249554 175710 249734 175798
rect 249842 175710 250022 175798
rect 250130 175710 250310 175798
rect 250564 175710 250744 175798
rect 360436 175710 360560 175798
rect 360814 175710 360994 175798
rect 361102 175710 361282 175798
rect 361390 175710 361570 175798
rect 361678 175710 361858 175798
rect 361966 175710 362146 175798
rect 362254 175710 362434 175798
rect 362542 175710 362722 175798
rect 362830 175710 363010 175798
rect 363264 175710 363444 175798
rect 363552 175710 363732 175798
rect 363840 175710 364020 175798
rect 364128 175710 364308 175798
rect 364416 175710 364596 175798
rect 364704 175710 364884 175798
rect 364992 175710 365172 175798
rect 365280 175710 365460 175798
rect 365714 175710 365894 175798
rect 366002 175710 366182 175798
rect 366290 175710 366470 175798
rect 366578 175710 366758 175798
rect 366866 175710 367046 175798
rect 367154 175710 367334 175798
rect 367442 175710 367622 175798
rect 367730 175710 367910 175798
rect 243214 175234 243394 175322
rect 243502 175234 243682 175322
rect 243790 175234 243970 175322
rect 244078 175234 244258 175322
rect 244366 175234 244546 175322
rect 244654 175234 244834 175322
rect 244942 175234 245122 175322
rect 245230 175234 245410 175322
rect 245664 175234 245844 175322
rect 245952 175234 246132 175322
rect 246240 175234 246420 175322
rect 246528 175234 246708 175322
rect 246816 175234 246996 175322
rect 247104 175234 247284 175322
rect 247392 175234 247572 175322
rect 247680 175234 247860 175322
rect 248114 175234 248294 175322
rect 248402 175234 248582 175322
rect 248690 175234 248870 175322
rect 248978 175234 249158 175322
rect 249266 175234 249446 175322
rect 249554 175234 249734 175322
rect 249842 175234 250022 175322
rect 250130 175234 250310 175322
rect 250564 175234 250744 175322
rect 360436 175234 360560 175322
rect 360814 175234 360994 175322
rect 361102 175234 361282 175322
rect 361390 175234 361570 175322
rect 361678 175234 361858 175322
rect 361966 175234 362146 175322
rect 362254 175234 362434 175322
rect 362542 175234 362722 175322
rect 362830 175234 363010 175322
rect 363264 175234 363444 175322
rect 363552 175234 363732 175322
rect 363840 175234 364020 175322
rect 364128 175234 364308 175322
rect 364416 175234 364596 175322
rect 364704 175234 364884 175322
rect 364992 175234 365172 175322
rect 365280 175234 365460 175322
rect 365714 175234 365894 175322
rect 366002 175234 366182 175322
rect 366290 175234 366470 175322
rect 366578 175234 366758 175322
rect 366866 175234 367046 175322
rect 367154 175234 367334 175322
rect 367442 175234 367622 175322
rect 367730 175234 367910 175322
rect 243214 175018 243394 175106
rect 243502 175018 243682 175106
rect 243790 175018 243970 175106
rect 244078 175018 244258 175106
rect 244366 175018 244546 175106
rect 244654 175018 244834 175106
rect 244942 175018 245122 175106
rect 245230 175018 245410 175106
rect 245664 175018 245844 175106
rect 245952 175018 246132 175106
rect 246240 175018 246420 175106
rect 246528 175018 246708 175106
rect 246816 175018 246996 175106
rect 247104 175018 247284 175106
rect 247392 175018 247572 175106
rect 247680 175018 247860 175106
rect 248114 175018 248294 175106
rect 248402 175018 248582 175106
rect 248690 175018 248870 175106
rect 248978 175018 249158 175106
rect 249266 175018 249446 175106
rect 249554 175018 249734 175106
rect 249842 175018 250022 175106
rect 250130 175018 250310 175106
rect 250564 175018 250744 175106
rect 360436 175018 360560 175106
rect 360814 175018 360994 175106
rect 361102 175018 361282 175106
rect 361390 175018 361570 175106
rect 361678 175018 361858 175106
rect 361966 175018 362146 175106
rect 362254 175018 362434 175106
rect 362542 175018 362722 175106
rect 362830 175018 363010 175106
rect 363264 175018 363444 175106
rect 363552 175018 363732 175106
rect 363840 175018 364020 175106
rect 364128 175018 364308 175106
rect 364416 175018 364596 175106
rect 364704 175018 364884 175106
rect 364992 175018 365172 175106
rect 365280 175018 365460 175106
rect 365714 175018 365894 175106
rect 366002 175018 366182 175106
rect 366290 175018 366470 175106
rect 366578 175018 366758 175106
rect 366866 175018 367046 175106
rect 367154 175018 367334 175106
rect 367442 175018 367622 175106
rect 367730 175018 367910 175106
rect 243214 174542 243394 174630
rect 243502 174542 243682 174630
rect 243790 174542 243970 174630
rect 244078 174542 244258 174630
rect 244366 174542 244546 174630
rect 244654 174542 244834 174630
rect 244942 174542 245122 174630
rect 245230 174542 245410 174630
rect 245664 174542 245844 174630
rect 245952 174542 246132 174630
rect 246240 174542 246420 174630
rect 246528 174542 246708 174630
rect 246816 174542 246996 174630
rect 247104 174542 247284 174630
rect 247392 174542 247572 174630
rect 247680 174542 247860 174630
rect 248114 174542 248294 174630
rect 248402 174542 248582 174630
rect 248690 174542 248870 174630
rect 248978 174542 249158 174630
rect 249266 174542 249446 174630
rect 249554 174542 249734 174630
rect 249842 174542 250022 174630
rect 250130 174542 250310 174630
rect 250564 174542 250744 174630
rect 360436 174542 360560 174630
rect 360814 174542 360994 174630
rect 361102 174542 361282 174630
rect 361390 174542 361570 174630
rect 361678 174542 361858 174630
rect 361966 174542 362146 174630
rect 362254 174542 362434 174630
rect 362542 174542 362722 174630
rect 362830 174542 363010 174630
rect 363264 174542 363444 174630
rect 363552 174542 363732 174630
rect 363840 174542 364020 174630
rect 364128 174542 364308 174630
rect 364416 174542 364596 174630
rect 364704 174542 364884 174630
rect 364992 174542 365172 174630
rect 365280 174542 365460 174630
rect 365714 174542 365894 174630
rect 366002 174542 366182 174630
rect 366290 174542 366470 174630
rect 366578 174542 366758 174630
rect 366866 174542 367046 174630
rect 367154 174542 367334 174630
rect 367442 174542 367622 174630
rect 367730 174542 367910 174630
rect 243214 174326 243394 174414
rect 243502 174326 243682 174414
rect 243790 174326 243970 174414
rect 244078 174326 244258 174414
rect 244366 174326 244546 174414
rect 244654 174326 244834 174414
rect 244942 174326 245122 174414
rect 245230 174326 245410 174414
rect 245664 174326 245844 174414
rect 245952 174326 246132 174414
rect 246240 174326 246420 174414
rect 246528 174326 246708 174414
rect 246816 174326 246996 174414
rect 247104 174326 247284 174414
rect 247392 174326 247572 174414
rect 247680 174326 247860 174414
rect 248114 174326 248294 174414
rect 248402 174326 248582 174414
rect 248690 174326 248870 174414
rect 248978 174326 249158 174414
rect 249266 174326 249446 174414
rect 249554 174326 249734 174414
rect 249842 174326 250022 174414
rect 250130 174326 250310 174414
rect 250564 174326 250744 174414
rect 360436 174326 360560 174414
rect 360814 174326 360994 174414
rect 361102 174326 361282 174414
rect 361390 174326 361570 174414
rect 361678 174326 361858 174414
rect 361966 174326 362146 174414
rect 362254 174326 362434 174414
rect 362542 174326 362722 174414
rect 362830 174326 363010 174414
rect 363264 174326 363444 174414
rect 363552 174326 363732 174414
rect 363840 174326 364020 174414
rect 364128 174326 364308 174414
rect 364416 174326 364596 174414
rect 364704 174326 364884 174414
rect 364992 174326 365172 174414
rect 365280 174326 365460 174414
rect 365714 174326 365894 174414
rect 366002 174326 366182 174414
rect 366290 174326 366470 174414
rect 366578 174326 366758 174414
rect 366866 174326 367046 174414
rect 367154 174326 367334 174414
rect 367442 174326 367622 174414
rect 367730 174326 367910 174414
rect 243214 173850 243394 173938
rect 243502 173850 243682 173938
rect 243790 173850 243970 173938
rect 244078 173850 244258 173938
rect 244366 173850 244546 173938
rect 244654 173850 244834 173938
rect 244942 173850 245122 173938
rect 245230 173850 245410 173938
rect 245664 173850 245844 173938
rect 245952 173850 246132 173938
rect 246240 173850 246420 173938
rect 246528 173850 246708 173938
rect 246816 173850 246996 173938
rect 247104 173850 247284 173938
rect 247392 173850 247572 173938
rect 247680 173850 247860 173938
rect 248114 173850 248294 173938
rect 248402 173850 248582 173938
rect 248690 173850 248870 173938
rect 248978 173850 249158 173938
rect 249266 173850 249446 173938
rect 249554 173850 249734 173938
rect 249842 173850 250022 173938
rect 250130 173850 250310 173938
rect 250564 173850 250744 173938
rect 360436 173850 360560 173938
rect 360814 173850 360994 173938
rect 361102 173850 361282 173938
rect 361390 173850 361570 173938
rect 361678 173850 361858 173938
rect 361966 173850 362146 173938
rect 362254 173850 362434 173938
rect 362542 173850 362722 173938
rect 362830 173850 363010 173938
rect 363264 173850 363444 173938
rect 363552 173850 363732 173938
rect 363840 173850 364020 173938
rect 364128 173850 364308 173938
rect 364416 173850 364596 173938
rect 364704 173850 364884 173938
rect 364992 173850 365172 173938
rect 365280 173850 365460 173938
rect 365714 173850 365894 173938
rect 366002 173850 366182 173938
rect 366290 173850 366470 173938
rect 366578 173850 366758 173938
rect 366866 173850 367046 173938
rect 367154 173850 367334 173938
rect 367442 173850 367622 173938
rect 367730 173850 367910 173938
rect 243214 173634 243394 173722
rect 243502 173634 243682 173722
rect 243790 173634 243970 173722
rect 244078 173634 244258 173722
rect 244366 173634 244546 173722
rect 244654 173634 244834 173722
rect 244942 173634 245122 173722
rect 245230 173634 245410 173722
rect 245664 173634 245844 173722
rect 245952 173634 246132 173722
rect 246240 173634 246420 173722
rect 246528 173634 246708 173722
rect 246816 173634 246996 173722
rect 247104 173634 247284 173722
rect 247392 173634 247572 173722
rect 247680 173634 247860 173722
rect 248114 173634 248294 173722
rect 248402 173634 248582 173722
rect 248690 173634 248870 173722
rect 248978 173634 249158 173722
rect 249266 173634 249446 173722
rect 249554 173634 249734 173722
rect 249842 173634 250022 173722
rect 250130 173634 250310 173722
rect 250564 173634 250744 173722
rect 360436 173634 360560 173722
rect 360814 173634 360994 173722
rect 361102 173634 361282 173722
rect 361390 173634 361570 173722
rect 361678 173634 361858 173722
rect 361966 173634 362146 173722
rect 362254 173634 362434 173722
rect 362542 173634 362722 173722
rect 362830 173634 363010 173722
rect 363264 173634 363444 173722
rect 363552 173634 363732 173722
rect 363840 173634 364020 173722
rect 364128 173634 364308 173722
rect 364416 173634 364596 173722
rect 364704 173634 364884 173722
rect 364992 173634 365172 173722
rect 365280 173634 365460 173722
rect 365714 173634 365894 173722
rect 366002 173634 366182 173722
rect 366290 173634 366470 173722
rect 366578 173634 366758 173722
rect 366866 173634 367046 173722
rect 367154 173634 367334 173722
rect 367442 173634 367622 173722
rect 367730 173634 367910 173722
rect 243214 173158 243394 173246
rect 243502 173158 243682 173246
rect 243790 173158 243970 173246
rect 244078 173158 244258 173246
rect 244366 173158 244546 173246
rect 244654 173158 244834 173246
rect 244942 173158 245122 173246
rect 245230 173158 245410 173246
rect 245664 173158 245844 173246
rect 245952 173158 246132 173246
rect 246240 173158 246420 173246
rect 246528 173158 246708 173246
rect 246816 173158 246996 173246
rect 247104 173158 247284 173246
rect 247392 173158 247572 173246
rect 247680 173158 247860 173246
rect 248114 173158 248294 173246
rect 248402 173158 248582 173246
rect 248690 173158 248870 173246
rect 248978 173158 249158 173246
rect 249266 173158 249446 173246
rect 249554 173158 249734 173246
rect 249842 173158 250022 173246
rect 250130 173158 250310 173246
rect 250564 173158 250744 173246
rect 360436 173158 360560 173246
rect 360814 173158 360994 173246
rect 361102 173158 361282 173246
rect 361390 173158 361570 173246
rect 361678 173158 361858 173246
rect 361966 173158 362146 173246
rect 362254 173158 362434 173246
rect 362542 173158 362722 173246
rect 362830 173158 363010 173246
rect 363264 173158 363444 173246
rect 363552 173158 363732 173246
rect 363840 173158 364020 173246
rect 364128 173158 364308 173246
rect 364416 173158 364596 173246
rect 364704 173158 364884 173246
rect 364992 173158 365172 173246
rect 365280 173158 365460 173246
rect 365714 173158 365894 173246
rect 366002 173158 366182 173246
rect 366290 173158 366470 173246
rect 366578 173158 366758 173246
rect 366866 173158 367046 173246
rect 367154 173158 367334 173246
rect 367442 173158 367622 173246
rect 367730 173158 367910 173246
rect 243214 172684 243394 172772
rect 243502 172684 243682 172772
rect 243790 172684 243970 172772
rect 244078 172684 244258 172772
rect 244366 172684 244546 172772
rect 244654 172684 244834 172772
rect 244942 172684 245122 172772
rect 245230 172684 245410 172772
rect 245664 172684 245844 172772
rect 245952 172684 246132 172772
rect 246240 172684 246420 172772
rect 246528 172684 246708 172772
rect 246816 172684 246996 172772
rect 247104 172684 247284 172772
rect 247392 172684 247572 172772
rect 247680 172684 247860 172772
rect 248114 172684 248294 172772
rect 248402 172684 248582 172772
rect 248690 172684 248870 172772
rect 248978 172684 249158 172772
rect 249266 172684 249446 172772
rect 249554 172684 249734 172772
rect 249842 172684 250022 172772
rect 250130 172684 250310 172772
rect 250564 172684 250744 172772
rect 360436 172684 360560 172772
rect 360814 172684 360994 172772
rect 361102 172684 361282 172772
rect 361390 172684 361570 172772
rect 361678 172684 361858 172772
rect 361966 172684 362146 172772
rect 362254 172684 362434 172772
rect 362542 172684 362722 172772
rect 362830 172684 363010 172772
rect 363264 172684 363444 172772
rect 363552 172684 363732 172772
rect 363840 172684 364020 172772
rect 364128 172684 364308 172772
rect 364416 172684 364596 172772
rect 364704 172684 364884 172772
rect 364992 172684 365172 172772
rect 365280 172684 365460 172772
rect 365714 172684 365894 172772
rect 366002 172684 366182 172772
rect 366290 172684 366470 172772
rect 366578 172684 366758 172772
rect 366866 172684 367046 172772
rect 367154 172684 367334 172772
rect 367442 172684 367622 172772
rect 367730 172684 367910 172772
rect 243214 172208 243394 172296
rect 243502 172208 243682 172296
rect 243790 172208 243970 172296
rect 244078 172208 244258 172296
rect 244366 172208 244546 172296
rect 244654 172208 244834 172296
rect 244942 172208 245122 172296
rect 245230 172208 245410 172296
rect 245664 172208 245844 172296
rect 245952 172208 246132 172296
rect 246240 172208 246420 172296
rect 246528 172208 246708 172296
rect 246816 172208 246996 172296
rect 247104 172208 247284 172296
rect 247392 172208 247572 172296
rect 247680 172208 247860 172296
rect 248114 172208 248294 172296
rect 248402 172208 248582 172296
rect 248690 172208 248870 172296
rect 248978 172208 249158 172296
rect 249266 172208 249446 172296
rect 249554 172208 249734 172296
rect 249842 172208 250022 172296
rect 250130 172208 250310 172296
rect 250564 172208 250744 172296
rect 360436 172208 360560 172296
rect 360814 172208 360994 172296
rect 361102 172208 361282 172296
rect 361390 172208 361570 172296
rect 361678 172208 361858 172296
rect 361966 172208 362146 172296
rect 362254 172208 362434 172296
rect 362542 172208 362722 172296
rect 362830 172208 363010 172296
rect 363264 172208 363444 172296
rect 363552 172208 363732 172296
rect 363840 172208 364020 172296
rect 364128 172208 364308 172296
rect 364416 172208 364596 172296
rect 364704 172208 364884 172296
rect 364992 172208 365172 172296
rect 365280 172208 365460 172296
rect 365714 172208 365894 172296
rect 366002 172208 366182 172296
rect 366290 172208 366470 172296
rect 366578 172208 366758 172296
rect 366866 172208 367046 172296
rect 367154 172208 367334 172296
rect 367442 172208 367622 172296
rect 367730 172208 367910 172296
rect 243214 171992 243394 172080
rect 243502 171992 243682 172080
rect 243790 171992 243970 172080
rect 244078 171992 244258 172080
rect 244366 171992 244546 172080
rect 244654 171992 244834 172080
rect 244942 171992 245122 172080
rect 245230 171992 245410 172080
rect 245664 171992 245844 172080
rect 245952 171992 246132 172080
rect 246240 171992 246420 172080
rect 246528 171992 246708 172080
rect 246816 171992 246996 172080
rect 247104 171992 247284 172080
rect 247392 171992 247572 172080
rect 247680 171992 247860 172080
rect 248114 171992 248294 172080
rect 248402 171992 248582 172080
rect 248690 171992 248870 172080
rect 248978 171992 249158 172080
rect 249266 171992 249446 172080
rect 249554 171992 249734 172080
rect 249842 171992 250022 172080
rect 250130 171992 250310 172080
rect 250564 171992 250744 172080
rect 360436 171992 360560 172080
rect 360814 171992 360994 172080
rect 361102 171992 361282 172080
rect 361390 171992 361570 172080
rect 361678 171992 361858 172080
rect 361966 171992 362146 172080
rect 362254 171992 362434 172080
rect 362542 171992 362722 172080
rect 362830 171992 363010 172080
rect 363264 171992 363444 172080
rect 363552 171992 363732 172080
rect 363840 171992 364020 172080
rect 364128 171992 364308 172080
rect 364416 171992 364596 172080
rect 364704 171992 364884 172080
rect 364992 171992 365172 172080
rect 365280 171992 365460 172080
rect 365714 171992 365894 172080
rect 366002 171992 366182 172080
rect 366290 171992 366470 172080
rect 366578 171992 366758 172080
rect 366866 171992 367046 172080
rect 367154 171992 367334 172080
rect 367442 171992 367622 172080
rect 367730 171992 367910 172080
rect 243214 171516 243394 171604
rect 243502 171516 243682 171604
rect 243790 171516 243970 171604
rect 244078 171516 244258 171604
rect 244366 171516 244546 171604
rect 244654 171516 244834 171604
rect 244942 171516 245122 171604
rect 245230 171516 245410 171604
rect 245664 171516 245844 171604
rect 245952 171516 246132 171604
rect 246240 171516 246420 171604
rect 246528 171516 246708 171604
rect 246816 171516 246996 171604
rect 247104 171516 247284 171604
rect 247392 171516 247572 171604
rect 247680 171516 247860 171604
rect 248114 171516 248294 171604
rect 248402 171516 248582 171604
rect 248690 171516 248870 171604
rect 248978 171516 249158 171604
rect 249266 171516 249446 171604
rect 249554 171516 249734 171604
rect 249842 171516 250022 171604
rect 250130 171516 250310 171604
rect 250564 171516 250744 171604
rect 360436 171516 360560 171604
rect 360814 171516 360994 171604
rect 361102 171516 361282 171604
rect 361390 171516 361570 171604
rect 361678 171516 361858 171604
rect 361966 171516 362146 171604
rect 362254 171516 362434 171604
rect 362542 171516 362722 171604
rect 362830 171516 363010 171604
rect 363264 171516 363444 171604
rect 363552 171516 363732 171604
rect 363840 171516 364020 171604
rect 364128 171516 364308 171604
rect 364416 171516 364596 171604
rect 364704 171516 364884 171604
rect 364992 171516 365172 171604
rect 365280 171516 365460 171604
rect 365714 171516 365894 171604
rect 366002 171516 366182 171604
rect 366290 171516 366470 171604
rect 366578 171516 366758 171604
rect 366866 171516 367046 171604
rect 367154 171516 367334 171604
rect 367442 171516 367622 171604
rect 367730 171516 367910 171604
rect 243214 171300 243394 171388
rect 243502 171300 243682 171388
rect 243790 171300 243970 171388
rect 244078 171300 244258 171388
rect 244366 171300 244546 171388
rect 244654 171300 244834 171388
rect 244942 171300 245122 171388
rect 245230 171300 245410 171388
rect 245664 171300 245844 171388
rect 245952 171300 246132 171388
rect 246240 171300 246420 171388
rect 246528 171300 246708 171388
rect 246816 171300 246996 171388
rect 247104 171300 247284 171388
rect 247392 171300 247572 171388
rect 247680 171300 247860 171388
rect 248114 171300 248294 171388
rect 248402 171300 248582 171388
rect 248690 171300 248870 171388
rect 248978 171300 249158 171388
rect 249266 171300 249446 171388
rect 249554 171300 249734 171388
rect 249842 171300 250022 171388
rect 250130 171300 250310 171388
rect 250564 171300 250744 171388
rect 360436 171300 360560 171388
rect 360814 171300 360994 171388
rect 361102 171300 361282 171388
rect 361390 171300 361570 171388
rect 361678 171300 361858 171388
rect 361966 171300 362146 171388
rect 362254 171300 362434 171388
rect 362542 171300 362722 171388
rect 362830 171300 363010 171388
rect 363264 171300 363444 171388
rect 363552 171300 363732 171388
rect 363840 171300 364020 171388
rect 364128 171300 364308 171388
rect 364416 171300 364596 171388
rect 364704 171300 364884 171388
rect 364992 171300 365172 171388
rect 365280 171300 365460 171388
rect 365714 171300 365894 171388
rect 366002 171300 366182 171388
rect 366290 171300 366470 171388
rect 366578 171300 366758 171388
rect 366866 171300 367046 171388
rect 367154 171300 367334 171388
rect 367442 171300 367622 171388
rect 367730 171300 367910 171388
rect 243214 170824 243394 170912
rect 243502 170824 243682 170912
rect 243790 170824 243970 170912
rect 244078 170824 244258 170912
rect 244366 170824 244546 170912
rect 244654 170824 244834 170912
rect 244942 170824 245122 170912
rect 245230 170824 245410 170912
rect 245664 170824 245844 170912
rect 245952 170824 246132 170912
rect 246240 170824 246420 170912
rect 246528 170824 246708 170912
rect 246816 170824 246996 170912
rect 247104 170824 247284 170912
rect 247392 170824 247572 170912
rect 247680 170824 247860 170912
rect 248114 170824 248294 170912
rect 248402 170824 248582 170912
rect 248690 170824 248870 170912
rect 248978 170824 249158 170912
rect 249266 170824 249446 170912
rect 249554 170824 249734 170912
rect 249842 170824 250022 170912
rect 250130 170824 250310 170912
rect 250564 170824 250744 170912
rect 360436 170824 360560 170912
rect 360814 170824 360994 170912
rect 361102 170824 361282 170912
rect 361390 170824 361570 170912
rect 361678 170824 361858 170912
rect 361966 170824 362146 170912
rect 362254 170824 362434 170912
rect 362542 170824 362722 170912
rect 362830 170824 363010 170912
rect 363264 170824 363444 170912
rect 363552 170824 363732 170912
rect 363840 170824 364020 170912
rect 364128 170824 364308 170912
rect 364416 170824 364596 170912
rect 364704 170824 364884 170912
rect 364992 170824 365172 170912
rect 365280 170824 365460 170912
rect 365714 170824 365894 170912
rect 366002 170824 366182 170912
rect 366290 170824 366470 170912
rect 366578 170824 366758 170912
rect 366866 170824 367046 170912
rect 367154 170824 367334 170912
rect 367442 170824 367622 170912
rect 367730 170824 367910 170912
rect 243214 170608 243394 170696
rect 243502 170608 243682 170696
rect 243790 170608 243970 170696
rect 244078 170608 244258 170696
rect 244366 170608 244546 170696
rect 244654 170608 244834 170696
rect 244942 170608 245122 170696
rect 245230 170608 245410 170696
rect 245664 170608 245844 170696
rect 245952 170608 246132 170696
rect 246240 170608 246420 170696
rect 246528 170608 246708 170696
rect 246816 170608 246996 170696
rect 247104 170608 247284 170696
rect 247392 170608 247572 170696
rect 247680 170608 247860 170696
rect 248114 170608 248294 170696
rect 248402 170608 248582 170696
rect 248690 170608 248870 170696
rect 248978 170608 249158 170696
rect 249266 170608 249446 170696
rect 249554 170608 249734 170696
rect 249842 170608 250022 170696
rect 250130 170608 250310 170696
rect 250564 170608 250744 170696
rect 360436 170608 360560 170696
rect 360814 170608 360994 170696
rect 361102 170608 361282 170696
rect 361390 170608 361570 170696
rect 361678 170608 361858 170696
rect 361966 170608 362146 170696
rect 362254 170608 362434 170696
rect 362542 170608 362722 170696
rect 362830 170608 363010 170696
rect 363264 170608 363444 170696
rect 363552 170608 363732 170696
rect 363840 170608 364020 170696
rect 364128 170608 364308 170696
rect 364416 170608 364596 170696
rect 364704 170608 364884 170696
rect 364992 170608 365172 170696
rect 365280 170608 365460 170696
rect 365714 170608 365894 170696
rect 366002 170608 366182 170696
rect 366290 170608 366470 170696
rect 366578 170608 366758 170696
rect 366866 170608 367046 170696
rect 367154 170608 367334 170696
rect 367442 170608 367622 170696
rect 367730 170608 367910 170696
rect 243214 170132 243394 170220
rect 243502 170132 243682 170220
rect 243790 170132 243970 170220
rect 244078 170132 244258 170220
rect 244366 170132 244546 170220
rect 244654 170132 244834 170220
rect 244942 170132 245122 170220
rect 245230 170132 245410 170220
rect 245664 170132 245844 170220
rect 245952 170132 246132 170220
rect 246240 170132 246420 170220
rect 246528 170132 246708 170220
rect 246816 170132 246996 170220
rect 247104 170132 247284 170220
rect 247392 170132 247572 170220
rect 247680 170132 247860 170220
rect 248114 170132 248294 170220
rect 248402 170132 248582 170220
rect 248690 170132 248870 170220
rect 248978 170132 249158 170220
rect 249266 170132 249446 170220
rect 249554 170132 249734 170220
rect 249842 170132 250022 170220
rect 250130 170132 250310 170220
rect 250564 170132 250744 170220
rect 360436 170132 360560 170220
rect 360814 170132 360994 170220
rect 361102 170132 361282 170220
rect 361390 170132 361570 170220
rect 361678 170132 361858 170220
rect 361966 170132 362146 170220
rect 362254 170132 362434 170220
rect 362542 170132 362722 170220
rect 362830 170132 363010 170220
rect 363264 170132 363444 170220
rect 363552 170132 363732 170220
rect 363840 170132 364020 170220
rect 364128 170132 364308 170220
rect 364416 170132 364596 170220
rect 364704 170132 364884 170220
rect 364992 170132 365172 170220
rect 365280 170132 365460 170220
rect 365714 170132 365894 170220
rect 366002 170132 366182 170220
rect 366290 170132 366470 170220
rect 366578 170132 366758 170220
rect 366866 170132 367046 170220
rect 367154 170132 367334 170220
rect 367442 170132 367622 170220
rect 367730 170132 367910 170220
rect 243214 169658 243394 169746
rect 243502 169658 243682 169746
rect 243790 169658 243970 169746
rect 244078 169658 244258 169746
rect 244366 169658 244546 169746
rect 244654 169658 244834 169746
rect 244942 169658 245122 169746
rect 245230 169658 245410 169746
rect 245664 169658 245844 169746
rect 245952 169658 246132 169746
rect 246240 169658 246420 169746
rect 246528 169658 246708 169746
rect 246816 169658 246996 169746
rect 247104 169658 247284 169746
rect 247392 169658 247572 169746
rect 247680 169658 247860 169746
rect 248114 169658 248294 169746
rect 248402 169658 248582 169746
rect 248690 169658 248870 169746
rect 248978 169658 249158 169746
rect 249266 169658 249446 169746
rect 249554 169658 249734 169746
rect 249842 169658 250022 169746
rect 250130 169658 250310 169746
rect 250564 169658 250744 169746
rect 360436 169658 360560 169746
rect 360814 169658 360994 169746
rect 361102 169658 361282 169746
rect 361390 169658 361570 169746
rect 361678 169658 361858 169746
rect 361966 169658 362146 169746
rect 362254 169658 362434 169746
rect 362542 169658 362722 169746
rect 362830 169658 363010 169746
rect 363264 169658 363444 169746
rect 363552 169658 363732 169746
rect 363840 169658 364020 169746
rect 364128 169658 364308 169746
rect 364416 169658 364596 169746
rect 364704 169658 364884 169746
rect 364992 169658 365172 169746
rect 365280 169658 365460 169746
rect 365714 169658 365894 169746
rect 366002 169658 366182 169746
rect 366290 169658 366470 169746
rect 366578 169658 366758 169746
rect 366866 169658 367046 169746
rect 367154 169658 367334 169746
rect 367442 169658 367622 169746
rect 367730 169658 367910 169746
rect 243214 169182 243394 169270
rect 243502 169182 243682 169270
rect 243790 169182 243970 169270
rect 244078 169182 244258 169270
rect 244366 169182 244546 169270
rect 244654 169182 244834 169270
rect 244942 169182 245122 169270
rect 245230 169182 245410 169270
rect 245664 169182 245844 169270
rect 245952 169182 246132 169270
rect 246240 169182 246420 169270
rect 246528 169182 246708 169270
rect 246816 169182 246996 169270
rect 247104 169182 247284 169270
rect 247392 169182 247572 169270
rect 247680 169182 247860 169270
rect 248114 169182 248294 169270
rect 248402 169182 248582 169270
rect 248690 169182 248870 169270
rect 248978 169182 249158 169270
rect 249266 169182 249446 169270
rect 249554 169182 249734 169270
rect 249842 169182 250022 169270
rect 250130 169182 250310 169270
rect 250564 169182 250744 169270
rect 360436 169182 360560 169270
rect 360814 169182 360994 169270
rect 361102 169182 361282 169270
rect 361390 169182 361570 169270
rect 361678 169182 361858 169270
rect 361966 169182 362146 169270
rect 362254 169182 362434 169270
rect 362542 169182 362722 169270
rect 362830 169182 363010 169270
rect 363264 169182 363444 169270
rect 363552 169182 363732 169270
rect 363840 169182 364020 169270
rect 364128 169182 364308 169270
rect 364416 169182 364596 169270
rect 364704 169182 364884 169270
rect 364992 169182 365172 169270
rect 365280 169182 365460 169270
rect 365714 169182 365894 169270
rect 366002 169182 366182 169270
rect 366290 169182 366470 169270
rect 366578 169182 366758 169270
rect 366866 169182 367046 169270
rect 367154 169182 367334 169270
rect 367442 169182 367622 169270
rect 367730 169182 367910 169270
rect 243214 168966 243394 169054
rect 243502 168966 243682 169054
rect 243790 168966 243970 169054
rect 244078 168966 244258 169054
rect 244366 168966 244546 169054
rect 244654 168966 244834 169054
rect 244942 168966 245122 169054
rect 245230 168966 245410 169054
rect 245664 168966 245844 169054
rect 245952 168966 246132 169054
rect 246240 168966 246420 169054
rect 246528 168966 246708 169054
rect 246816 168966 246996 169054
rect 247104 168966 247284 169054
rect 247392 168966 247572 169054
rect 247680 168966 247860 169054
rect 248114 168966 248294 169054
rect 248402 168966 248582 169054
rect 248690 168966 248870 169054
rect 248978 168966 249158 169054
rect 249266 168966 249446 169054
rect 249554 168966 249734 169054
rect 249842 168966 250022 169054
rect 250130 168966 250310 169054
rect 250564 168966 250744 169054
rect 360436 168966 360560 169054
rect 360814 168966 360994 169054
rect 361102 168966 361282 169054
rect 361390 168966 361570 169054
rect 361678 168966 361858 169054
rect 361966 168966 362146 169054
rect 362254 168966 362434 169054
rect 362542 168966 362722 169054
rect 362830 168966 363010 169054
rect 363264 168966 363444 169054
rect 363552 168966 363732 169054
rect 363840 168966 364020 169054
rect 364128 168966 364308 169054
rect 364416 168966 364596 169054
rect 364704 168966 364884 169054
rect 364992 168966 365172 169054
rect 365280 168966 365460 169054
rect 365714 168966 365894 169054
rect 366002 168966 366182 169054
rect 366290 168966 366470 169054
rect 366578 168966 366758 169054
rect 366866 168966 367046 169054
rect 367154 168966 367334 169054
rect 367442 168966 367622 169054
rect 367730 168966 367910 169054
rect 243214 168490 243394 168578
rect 243502 168490 243682 168578
rect 243790 168490 243970 168578
rect 244078 168490 244258 168578
rect 244366 168490 244546 168578
rect 244654 168490 244834 168578
rect 244942 168490 245122 168578
rect 245230 168490 245410 168578
rect 245664 168490 245844 168578
rect 245952 168490 246132 168578
rect 246240 168490 246420 168578
rect 246528 168490 246708 168578
rect 246816 168490 246996 168578
rect 247104 168490 247284 168578
rect 247392 168490 247572 168578
rect 247680 168490 247860 168578
rect 248114 168490 248294 168578
rect 248402 168490 248582 168578
rect 248690 168490 248870 168578
rect 248978 168490 249158 168578
rect 249266 168490 249446 168578
rect 249554 168490 249734 168578
rect 249842 168490 250022 168578
rect 250130 168490 250310 168578
rect 250564 168490 250744 168578
rect 360436 168490 360560 168578
rect 360814 168490 360994 168578
rect 361102 168490 361282 168578
rect 361390 168490 361570 168578
rect 361678 168490 361858 168578
rect 361966 168490 362146 168578
rect 362254 168490 362434 168578
rect 362542 168490 362722 168578
rect 362830 168490 363010 168578
rect 363264 168490 363444 168578
rect 363552 168490 363732 168578
rect 363840 168490 364020 168578
rect 364128 168490 364308 168578
rect 364416 168490 364596 168578
rect 364704 168490 364884 168578
rect 364992 168490 365172 168578
rect 365280 168490 365460 168578
rect 365714 168490 365894 168578
rect 366002 168490 366182 168578
rect 366290 168490 366470 168578
rect 366578 168490 366758 168578
rect 366866 168490 367046 168578
rect 367154 168490 367334 168578
rect 367442 168490 367622 168578
rect 367730 168490 367910 168578
rect 243214 168274 243394 168362
rect 243502 168274 243682 168362
rect 243790 168274 243970 168362
rect 244078 168274 244258 168362
rect 244366 168274 244546 168362
rect 244654 168274 244834 168362
rect 244942 168274 245122 168362
rect 245230 168274 245410 168362
rect 245664 168274 245844 168362
rect 245952 168274 246132 168362
rect 246240 168274 246420 168362
rect 246528 168274 246708 168362
rect 246816 168274 246996 168362
rect 247104 168274 247284 168362
rect 247392 168274 247572 168362
rect 247680 168274 247860 168362
rect 248114 168274 248294 168362
rect 248402 168274 248582 168362
rect 248690 168274 248870 168362
rect 248978 168274 249158 168362
rect 249266 168274 249446 168362
rect 249554 168274 249734 168362
rect 249842 168274 250022 168362
rect 250130 168274 250310 168362
rect 250564 168274 250744 168362
rect 360436 168274 360560 168362
rect 360814 168274 360994 168362
rect 361102 168274 361282 168362
rect 361390 168274 361570 168362
rect 361678 168274 361858 168362
rect 361966 168274 362146 168362
rect 362254 168274 362434 168362
rect 362542 168274 362722 168362
rect 362830 168274 363010 168362
rect 363264 168274 363444 168362
rect 363552 168274 363732 168362
rect 363840 168274 364020 168362
rect 364128 168274 364308 168362
rect 364416 168274 364596 168362
rect 364704 168274 364884 168362
rect 364992 168274 365172 168362
rect 365280 168274 365460 168362
rect 365714 168274 365894 168362
rect 366002 168274 366182 168362
rect 366290 168274 366470 168362
rect 366578 168274 366758 168362
rect 366866 168274 367046 168362
rect 367154 168274 367334 168362
rect 367442 168274 367622 168362
rect 367730 168274 367910 168362
rect 243214 167798 243394 167886
rect 243502 167798 243682 167886
rect 243790 167798 243970 167886
rect 244078 167798 244258 167886
rect 244366 167798 244546 167886
rect 244654 167798 244834 167886
rect 244942 167798 245122 167886
rect 245230 167798 245410 167886
rect 245664 167798 245844 167886
rect 245952 167798 246132 167886
rect 246240 167798 246420 167886
rect 246528 167798 246708 167886
rect 246816 167798 246996 167886
rect 247104 167798 247284 167886
rect 247392 167798 247572 167886
rect 247680 167798 247860 167886
rect 248114 167798 248294 167886
rect 248402 167798 248582 167886
rect 248690 167798 248870 167886
rect 248978 167798 249158 167886
rect 249266 167798 249446 167886
rect 249554 167798 249734 167886
rect 249842 167798 250022 167886
rect 250130 167798 250310 167886
rect 250564 167798 250744 167886
rect 360436 167798 360560 167886
rect 360814 167798 360994 167886
rect 361102 167798 361282 167886
rect 361390 167798 361570 167886
rect 361678 167798 361858 167886
rect 361966 167798 362146 167886
rect 362254 167798 362434 167886
rect 362542 167798 362722 167886
rect 362830 167798 363010 167886
rect 363264 167798 363444 167886
rect 363552 167798 363732 167886
rect 363840 167798 364020 167886
rect 364128 167798 364308 167886
rect 364416 167798 364596 167886
rect 364704 167798 364884 167886
rect 364992 167798 365172 167886
rect 365280 167798 365460 167886
rect 365714 167798 365894 167886
rect 366002 167798 366182 167886
rect 366290 167798 366470 167886
rect 366578 167798 366758 167886
rect 366866 167798 367046 167886
rect 367154 167798 367334 167886
rect 367442 167798 367622 167886
rect 367730 167798 367910 167886
rect 243214 167582 243394 167670
rect 243502 167582 243682 167670
rect 243790 167582 243970 167670
rect 244078 167582 244258 167670
rect 244366 167582 244546 167670
rect 244654 167582 244834 167670
rect 244942 167582 245122 167670
rect 245230 167582 245410 167670
rect 245664 167582 245844 167670
rect 245952 167582 246132 167670
rect 246240 167582 246420 167670
rect 246528 167582 246708 167670
rect 246816 167582 246996 167670
rect 247104 167582 247284 167670
rect 247392 167582 247572 167670
rect 247680 167582 247860 167670
rect 248114 167582 248294 167670
rect 248402 167582 248582 167670
rect 248690 167582 248870 167670
rect 248978 167582 249158 167670
rect 249266 167582 249446 167670
rect 249554 167582 249734 167670
rect 249842 167582 250022 167670
rect 250130 167582 250310 167670
rect 250564 167582 250744 167670
rect 360436 167582 360560 167670
rect 360814 167582 360994 167670
rect 361102 167582 361282 167670
rect 361390 167582 361570 167670
rect 361678 167582 361858 167670
rect 361966 167582 362146 167670
rect 362254 167582 362434 167670
rect 362542 167582 362722 167670
rect 362830 167582 363010 167670
rect 363264 167582 363444 167670
rect 363552 167582 363732 167670
rect 363840 167582 364020 167670
rect 364128 167582 364308 167670
rect 364416 167582 364596 167670
rect 364704 167582 364884 167670
rect 364992 167582 365172 167670
rect 365280 167582 365460 167670
rect 365714 167582 365894 167670
rect 366002 167582 366182 167670
rect 366290 167582 366470 167670
rect 366578 167582 366758 167670
rect 366866 167582 367046 167670
rect 367154 167582 367334 167670
rect 367442 167582 367622 167670
rect 367730 167582 367910 167670
rect 243214 167106 243394 167194
rect 243502 167106 243682 167194
rect 243790 167106 243970 167194
rect 244078 167106 244258 167194
rect 244366 167106 244546 167194
rect 244654 167106 244834 167194
rect 244942 167106 245122 167194
rect 245230 167106 245410 167194
rect 245664 167106 245844 167194
rect 245952 167106 246132 167194
rect 246240 167106 246420 167194
rect 246528 167106 246708 167194
rect 246816 167106 246996 167194
rect 247104 167106 247284 167194
rect 247392 167106 247572 167194
rect 247680 167106 247860 167194
rect 248114 167106 248294 167194
rect 248402 167106 248582 167194
rect 248690 167106 248870 167194
rect 248978 167106 249158 167194
rect 249266 167106 249446 167194
rect 249554 167106 249734 167194
rect 249842 167106 250022 167194
rect 250130 167106 250310 167194
rect 250564 167106 250744 167194
rect 360436 167106 360560 167194
rect 360814 167106 360994 167194
rect 361102 167106 361282 167194
rect 361390 167106 361570 167194
rect 361678 167106 361858 167194
rect 361966 167106 362146 167194
rect 362254 167106 362434 167194
rect 362542 167106 362722 167194
rect 362830 167106 363010 167194
rect 363264 167106 363444 167194
rect 363552 167106 363732 167194
rect 363840 167106 364020 167194
rect 364128 167106 364308 167194
rect 364416 167106 364596 167194
rect 364704 167106 364884 167194
rect 364992 167106 365172 167194
rect 365280 167106 365460 167194
rect 365714 167106 365894 167194
rect 366002 167106 366182 167194
rect 366290 167106 366470 167194
rect 366578 167106 366758 167194
rect 366866 167106 367046 167194
rect 367154 167106 367334 167194
rect 367442 167106 367622 167194
rect 367730 167106 367910 167194
rect 243214 166632 243394 166720
rect 243502 166632 243682 166720
rect 243790 166632 243970 166720
rect 244078 166632 244258 166720
rect 244366 166632 244546 166720
rect 244654 166632 244834 166720
rect 244942 166632 245122 166720
rect 245230 166632 245410 166720
rect 245664 166632 245844 166720
rect 245952 166632 246132 166720
rect 246240 166632 246420 166720
rect 246528 166632 246708 166720
rect 246816 166632 246996 166720
rect 247104 166632 247284 166720
rect 247392 166632 247572 166720
rect 247680 166632 247860 166720
rect 248114 166632 248294 166720
rect 248402 166632 248582 166720
rect 248690 166632 248870 166720
rect 248978 166632 249158 166720
rect 249266 166632 249446 166720
rect 249554 166632 249734 166720
rect 249842 166632 250022 166720
rect 250130 166632 250310 166720
rect 250564 166632 250744 166720
rect 360436 166632 360560 166720
rect 360814 166632 360994 166720
rect 361102 166632 361282 166720
rect 361390 166632 361570 166720
rect 361678 166632 361858 166720
rect 361966 166632 362146 166720
rect 362254 166632 362434 166720
rect 362542 166632 362722 166720
rect 362830 166632 363010 166720
rect 363264 166632 363444 166720
rect 363552 166632 363732 166720
rect 363840 166632 364020 166720
rect 364128 166632 364308 166720
rect 364416 166632 364596 166720
rect 364704 166632 364884 166720
rect 364992 166632 365172 166720
rect 365280 166632 365460 166720
rect 365714 166632 365894 166720
rect 366002 166632 366182 166720
rect 366290 166632 366470 166720
rect 366578 166632 366758 166720
rect 366866 166632 367046 166720
rect 367154 166632 367334 166720
rect 367442 166632 367622 166720
rect 367730 166632 367910 166720
rect 243214 166156 243394 166244
rect 243502 166156 243682 166244
rect 243790 166156 243970 166244
rect 244078 166156 244258 166244
rect 244366 166156 244546 166244
rect 244654 166156 244834 166244
rect 244942 166156 245122 166244
rect 245230 166156 245410 166244
rect 245664 166156 245844 166244
rect 245952 166156 246132 166244
rect 246240 166156 246420 166244
rect 246528 166156 246708 166244
rect 246816 166156 246996 166244
rect 247104 166156 247284 166244
rect 247392 166156 247572 166244
rect 247680 166156 247860 166244
rect 248114 166156 248294 166244
rect 248402 166156 248582 166244
rect 248690 166156 248870 166244
rect 248978 166156 249158 166244
rect 249266 166156 249446 166244
rect 249554 166156 249734 166244
rect 249842 166156 250022 166244
rect 250130 166156 250310 166244
rect 250564 166156 250744 166244
rect 360436 166156 360560 166244
rect 360814 166156 360994 166244
rect 361102 166156 361282 166244
rect 361390 166156 361570 166244
rect 361678 166156 361858 166244
rect 361966 166156 362146 166244
rect 362254 166156 362434 166244
rect 362542 166156 362722 166244
rect 362830 166156 363010 166244
rect 363264 166156 363444 166244
rect 363552 166156 363732 166244
rect 363840 166156 364020 166244
rect 364128 166156 364308 166244
rect 364416 166156 364596 166244
rect 364704 166156 364884 166244
rect 364992 166156 365172 166244
rect 365280 166156 365460 166244
rect 365714 166156 365894 166244
rect 366002 166156 366182 166244
rect 366290 166156 366470 166244
rect 366578 166156 366758 166244
rect 366866 166156 367046 166244
rect 367154 166156 367334 166244
rect 367442 166156 367622 166244
rect 367730 166156 367910 166244
rect 243214 165940 243394 166028
rect 243502 165940 243682 166028
rect 243790 165940 243970 166028
rect 244078 165940 244258 166028
rect 244366 165940 244546 166028
rect 244654 165940 244834 166028
rect 244942 165940 245122 166028
rect 245230 165940 245410 166028
rect 245664 165940 245844 166028
rect 245952 165940 246132 166028
rect 246240 165940 246420 166028
rect 246528 165940 246708 166028
rect 246816 165940 246996 166028
rect 247104 165940 247284 166028
rect 247392 165940 247572 166028
rect 247680 165940 247860 166028
rect 248114 165940 248294 166028
rect 248402 165940 248582 166028
rect 248690 165940 248870 166028
rect 248978 165940 249158 166028
rect 249266 165940 249446 166028
rect 249554 165940 249734 166028
rect 249842 165940 250022 166028
rect 250130 165940 250310 166028
rect 250564 165940 250744 166028
rect 360436 165940 360560 166028
rect 360814 165940 360994 166028
rect 361102 165940 361282 166028
rect 361390 165940 361570 166028
rect 361678 165940 361858 166028
rect 361966 165940 362146 166028
rect 362254 165940 362434 166028
rect 362542 165940 362722 166028
rect 362830 165940 363010 166028
rect 363264 165940 363444 166028
rect 363552 165940 363732 166028
rect 363840 165940 364020 166028
rect 364128 165940 364308 166028
rect 364416 165940 364596 166028
rect 364704 165940 364884 166028
rect 364992 165940 365172 166028
rect 365280 165940 365460 166028
rect 365714 165940 365894 166028
rect 366002 165940 366182 166028
rect 366290 165940 366470 166028
rect 366578 165940 366758 166028
rect 366866 165940 367046 166028
rect 367154 165940 367334 166028
rect 367442 165940 367622 166028
rect 367730 165940 367910 166028
rect 243214 165464 243394 165552
rect 243502 165464 243682 165552
rect 243790 165464 243970 165552
rect 244078 165464 244258 165552
rect 244366 165464 244546 165552
rect 244654 165464 244834 165552
rect 244942 165464 245122 165552
rect 245230 165464 245410 165552
rect 245664 165464 245844 165552
rect 245952 165464 246132 165552
rect 246240 165464 246420 165552
rect 246528 165464 246708 165552
rect 246816 165464 246996 165552
rect 247104 165464 247284 165552
rect 247392 165464 247572 165552
rect 247680 165464 247860 165552
rect 248114 165464 248294 165552
rect 248402 165464 248582 165552
rect 248690 165464 248870 165552
rect 248978 165464 249158 165552
rect 249266 165464 249446 165552
rect 249554 165464 249734 165552
rect 249842 165464 250022 165552
rect 250130 165464 250310 165552
rect 250564 165464 250744 165552
rect 360436 165464 360560 165552
rect 360814 165464 360994 165552
rect 361102 165464 361282 165552
rect 361390 165464 361570 165552
rect 361678 165464 361858 165552
rect 361966 165464 362146 165552
rect 362254 165464 362434 165552
rect 362542 165464 362722 165552
rect 362830 165464 363010 165552
rect 363264 165464 363444 165552
rect 363552 165464 363732 165552
rect 363840 165464 364020 165552
rect 364128 165464 364308 165552
rect 364416 165464 364596 165552
rect 364704 165464 364884 165552
rect 364992 165464 365172 165552
rect 365280 165464 365460 165552
rect 365714 165464 365894 165552
rect 366002 165464 366182 165552
rect 366290 165464 366470 165552
rect 366578 165464 366758 165552
rect 366866 165464 367046 165552
rect 367154 165464 367334 165552
rect 367442 165464 367622 165552
rect 367730 165464 367910 165552
rect 243214 165248 243394 165336
rect 243502 165248 243682 165336
rect 243790 165248 243970 165336
rect 244078 165248 244258 165336
rect 244366 165248 244546 165336
rect 244654 165248 244834 165336
rect 244942 165248 245122 165336
rect 245230 165248 245410 165336
rect 245664 165248 245844 165336
rect 245952 165248 246132 165336
rect 246240 165248 246420 165336
rect 246528 165248 246708 165336
rect 246816 165248 246996 165336
rect 247104 165248 247284 165336
rect 247392 165248 247572 165336
rect 247680 165248 247860 165336
rect 248114 165248 248294 165336
rect 248402 165248 248582 165336
rect 248690 165248 248870 165336
rect 248978 165248 249158 165336
rect 249266 165248 249446 165336
rect 249554 165248 249734 165336
rect 249842 165248 250022 165336
rect 250130 165248 250310 165336
rect 250564 165248 250744 165336
rect 360436 165248 360560 165336
rect 360814 165248 360994 165336
rect 361102 165248 361282 165336
rect 361390 165248 361570 165336
rect 361678 165248 361858 165336
rect 361966 165248 362146 165336
rect 362254 165248 362434 165336
rect 362542 165248 362722 165336
rect 362830 165248 363010 165336
rect 363264 165248 363444 165336
rect 363552 165248 363732 165336
rect 363840 165248 364020 165336
rect 364128 165248 364308 165336
rect 364416 165248 364596 165336
rect 364704 165248 364884 165336
rect 364992 165248 365172 165336
rect 365280 165248 365460 165336
rect 365714 165248 365894 165336
rect 366002 165248 366182 165336
rect 366290 165248 366470 165336
rect 366578 165248 366758 165336
rect 366866 165248 367046 165336
rect 367154 165248 367334 165336
rect 367442 165248 367622 165336
rect 367730 165248 367910 165336
rect 243214 164772 243394 164860
rect 243502 164772 243682 164860
rect 243790 164772 243970 164860
rect 244078 164772 244258 164860
rect 244366 164772 244546 164860
rect 244654 164772 244834 164860
rect 244942 164772 245122 164860
rect 245230 164772 245410 164860
rect 245664 164772 245844 164860
rect 245952 164772 246132 164860
rect 246240 164772 246420 164860
rect 246528 164772 246708 164860
rect 246816 164772 246996 164860
rect 247104 164772 247284 164860
rect 247392 164772 247572 164860
rect 247680 164772 247860 164860
rect 248114 164772 248294 164860
rect 248402 164772 248582 164860
rect 248690 164772 248870 164860
rect 248978 164772 249158 164860
rect 249266 164772 249446 164860
rect 249554 164772 249734 164860
rect 249842 164772 250022 164860
rect 250130 164772 250310 164860
rect 250564 164772 250744 164860
rect 360436 164772 360560 164860
rect 360814 164772 360994 164860
rect 361102 164772 361282 164860
rect 361390 164772 361570 164860
rect 361678 164772 361858 164860
rect 361966 164772 362146 164860
rect 362254 164772 362434 164860
rect 362542 164772 362722 164860
rect 362830 164772 363010 164860
rect 363264 164772 363444 164860
rect 363552 164772 363732 164860
rect 363840 164772 364020 164860
rect 364128 164772 364308 164860
rect 364416 164772 364596 164860
rect 364704 164772 364884 164860
rect 364992 164772 365172 164860
rect 365280 164772 365460 164860
rect 365714 164772 365894 164860
rect 366002 164772 366182 164860
rect 366290 164772 366470 164860
rect 366578 164772 366758 164860
rect 366866 164772 367046 164860
rect 367154 164772 367334 164860
rect 367442 164772 367622 164860
rect 367730 164772 367910 164860
rect 243214 164556 243394 164644
rect 243502 164556 243682 164644
rect 243790 164556 243970 164644
rect 244078 164556 244258 164644
rect 244366 164556 244546 164644
rect 244654 164556 244834 164644
rect 244942 164556 245122 164644
rect 245230 164556 245410 164644
rect 245664 164556 245844 164644
rect 245952 164556 246132 164644
rect 246240 164556 246420 164644
rect 246528 164556 246708 164644
rect 246816 164556 246996 164644
rect 247104 164556 247284 164644
rect 247392 164556 247572 164644
rect 247680 164556 247860 164644
rect 248114 164556 248294 164644
rect 248402 164556 248582 164644
rect 248690 164556 248870 164644
rect 248978 164556 249158 164644
rect 249266 164556 249446 164644
rect 249554 164556 249734 164644
rect 249842 164556 250022 164644
rect 250130 164556 250310 164644
rect 250564 164556 250744 164644
rect 360436 164556 360560 164644
rect 360814 164556 360994 164644
rect 361102 164556 361282 164644
rect 361390 164556 361570 164644
rect 361678 164556 361858 164644
rect 361966 164556 362146 164644
rect 362254 164556 362434 164644
rect 362542 164556 362722 164644
rect 362830 164556 363010 164644
rect 363264 164556 363444 164644
rect 363552 164556 363732 164644
rect 363840 164556 364020 164644
rect 364128 164556 364308 164644
rect 364416 164556 364596 164644
rect 364704 164556 364884 164644
rect 364992 164556 365172 164644
rect 365280 164556 365460 164644
rect 365714 164556 365894 164644
rect 366002 164556 366182 164644
rect 366290 164556 366470 164644
rect 366578 164556 366758 164644
rect 366866 164556 367046 164644
rect 367154 164556 367334 164644
rect 367442 164556 367622 164644
rect 367730 164556 367910 164644
rect 243214 164080 243394 164168
rect 243502 164080 243682 164168
rect 243790 164080 243970 164168
rect 244078 164080 244258 164168
rect 244366 164080 244546 164168
rect 244654 164080 244834 164168
rect 244942 164080 245122 164168
rect 245230 164080 245410 164168
rect 245664 164080 245844 164168
rect 245952 164080 246132 164168
rect 246240 164080 246420 164168
rect 246528 164080 246708 164168
rect 246816 164080 246996 164168
rect 247104 164080 247284 164168
rect 247392 164080 247572 164168
rect 247680 164080 247860 164168
rect 248114 164080 248294 164168
rect 248402 164080 248582 164168
rect 248690 164080 248870 164168
rect 248978 164080 249158 164168
rect 249266 164080 249446 164168
rect 249554 164080 249734 164168
rect 249842 164080 250022 164168
rect 250130 164080 250310 164168
rect 250564 164080 250744 164168
rect 360436 164080 360560 164168
rect 360814 164080 360994 164168
rect 361102 164080 361282 164168
rect 361390 164080 361570 164168
rect 361678 164080 361858 164168
rect 361966 164080 362146 164168
rect 362254 164080 362434 164168
rect 362542 164080 362722 164168
rect 362830 164080 363010 164168
rect 363264 164080 363444 164168
rect 363552 164080 363732 164168
rect 363840 164080 364020 164168
rect 364128 164080 364308 164168
rect 364416 164080 364596 164168
rect 364704 164080 364884 164168
rect 364992 164080 365172 164168
rect 365280 164080 365460 164168
rect 365714 164080 365894 164168
rect 366002 164080 366182 164168
rect 366290 164080 366470 164168
rect 366578 164080 366758 164168
rect 366866 164080 367046 164168
rect 367154 164080 367334 164168
rect 367442 164080 367622 164168
rect 367730 164080 367910 164168
rect 243214 163606 243394 163694
rect 243502 163606 243682 163694
rect 243790 163606 243970 163694
rect 244078 163606 244258 163694
rect 244366 163606 244546 163694
rect 244654 163606 244834 163694
rect 244942 163606 245122 163694
rect 245230 163606 245410 163694
rect 245664 163606 245844 163694
rect 245952 163606 246132 163694
rect 246240 163606 246420 163694
rect 246528 163606 246708 163694
rect 246816 163606 246996 163694
rect 247104 163606 247284 163694
rect 247392 163606 247572 163694
rect 247680 163606 247860 163694
rect 248114 163606 248294 163694
rect 248402 163606 248582 163694
rect 248690 163606 248870 163694
rect 248978 163606 249158 163694
rect 249266 163606 249446 163694
rect 249554 163606 249734 163694
rect 249842 163606 250022 163694
rect 250130 163606 250310 163694
rect 250564 163606 250744 163694
rect 360436 163606 360560 163694
rect 360814 163606 360994 163694
rect 361102 163606 361282 163694
rect 361390 163606 361570 163694
rect 361678 163606 361858 163694
rect 361966 163606 362146 163694
rect 362254 163606 362434 163694
rect 362542 163606 362722 163694
rect 362830 163606 363010 163694
rect 363264 163606 363444 163694
rect 363552 163606 363732 163694
rect 363840 163606 364020 163694
rect 364128 163606 364308 163694
rect 364416 163606 364596 163694
rect 364704 163606 364884 163694
rect 364992 163606 365172 163694
rect 365280 163606 365460 163694
rect 365714 163606 365894 163694
rect 366002 163606 366182 163694
rect 366290 163606 366470 163694
rect 366578 163606 366758 163694
rect 366866 163606 367046 163694
rect 367154 163606 367334 163694
rect 367442 163606 367622 163694
rect 367730 163606 367910 163694
rect 243214 163130 243394 163218
rect 243502 163130 243682 163218
rect 243790 163130 243970 163218
rect 244078 163130 244258 163218
rect 244366 163130 244546 163218
rect 244654 163130 244834 163218
rect 244942 163130 245122 163218
rect 245230 163130 245410 163218
rect 245664 163130 245844 163218
rect 245952 163130 246132 163218
rect 246240 163130 246420 163218
rect 246528 163130 246708 163218
rect 246816 163130 246996 163218
rect 247104 163130 247284 163218
rect 247392 163130 247572 163218
rect 247680 163130 247860 163218
rect 248114 163130 248294 163218
rect 248402 163130 248582 163218
rect 248690 163130 248870 163218
rect 248978 163130 249158 163218
rect 249266 163130 249446 163218
rect 249554 163130 249734 163218
rect 249842 163130 250022 163218
rect 250130 163130 250310 163218
rect 250564 163130 250744 163218
rect 360436 163130 360560 163218
rect 360814 163130 360994 163218
rect 361102 163130 361282 163218
rect 361390 163130 361570 163218
rect 361678 163130 361858 163218
rect 361966 163130 362146 163218
rect 362254 163130 362434 163218
rect 362542 163130 362722 163218
rect 362830 163130 363010 163218
rect 363264 163130 363444 163218
rect 363552 163130 363732 163218
rect 363840 163130 364020 163218
rect 364128 163130 364308 163218
rect 364416 163130 364596 163218
rect 364704 163130 364884 163218
rect 364992 163130 365172 163218
rect 365280 163130 365460 163218
rect 365714 163130 365894 163218
rect 366002 163130 366182 163218
rect 366290 163130 366470 163218
rect 366578 163130 366758 163218
rect 366866 163130 367046 163218
rect 367154 163130 367334 163218
rect 367442 163130 367622 163218
rect 367730 163130 367910 163218
rect 243214 162914 243394 163002
rect 243502 162914 243682 163002
rect 243790 162914 243970 163002
rect 244078 162914 244258 163002
rect 244366 162914 244546 163002
rect 244654 162914 244834 163002
rect 244942 162914 245122 163002
rect 245230 162914 245410 163002
rect 245664 162914 245844 163002
rect 245952 162914 246132 163002
rect 246240 162914 246420 163002
rect 246528 162914 246708 163002
rect 246816 162914 246996 163002
rect 247104 162914 247284 163002
rect 247392 162914 247572 163002
rect 247680 162914 247860 163002
rect 248114 162914 248294 163002
rect 248402 162914 248582 163002
rect 248690 162914 248870 163002
rect 248978 162914 249158 163002
rect 249266 162914 249446 163002
rect 249554 162914 249734 163002
rect 249842 162914 250022 163002
rect 250130 162914 250310 163002
rect 250564 162914 250744 163002
rect 360436 162914 360560 163002
rect 360814 162914 360994 163002
rect 361102 162914 361282 163002
rect 361390 162914 361570 163002
rect 361678 162914 361858 163002
rect 361966 162914 362146 163002
rect 362254 162914 362434 163002
rect 362542 162914 362722 163002
rect 362830 162914 363010 163002
rect 363264 162914 363444 163002
rect 363552 162914 363732 163002
rect 363840 162914 364020 163002
rect 364128 162914 364308 163002
rect 364416 162914 364596 163002
rect 364704 162914 364884 163002
rect 364992 162914 365172 163002
rect 365280 162914 365460 163002
rect 365714 162914 365894 163002
rect 366002 162914 366182 163002
rect 366290 162914 366470 163002
rect 366578 162914 366758 163002
rect 366866 162914 367046 163002
rect 367154 162914 367334 163002
rect 367442 162914 367622 163002
rect 367730 162914 367910 163002
rect 243214 162438 243394 162526
rect 243502 162438 243682 162526
rect 243790 162438 243970 162526
rect 244078 162438 244258 162526
rect 244366 162438 244546 162526
rect 244654 162438 244834 162526
rect 244942 162438 245122 162526
rect 245230 162438 245410 162526
rect 245664 162438 245844 162526
rect 245952 162438 246132 162526
rect 246240 162438 246420 162526
rect 246528 162438 246708 162526
rect 246816 162438 246996 162526
rect 247104 162438 247284 162526
rect 247392 162438 247572 162526
rect 247680 162438 247860 162526
rect 248114 162438 248294 162526
rect 248402 162438 248582 162526
rect 248690 162438 248870 162526
rect 248978 162438 249158 162526
rect 249266 162438 249446 162526
rect 249554 162438 249734 162526
rect 249842 162438 250022 162526
rect 250130 162438 250310 162526
rect 250564 162438 250744 162526
rect 360436 162438 360560 162526
rect 360814 162438 360994 162526
rect 361102 162438 361282 162526
rect 361390 162438 361570 162526
rect 361678 162438 361858 162526
rect 361966 162438 362146 162526
rect 362254 162438 362434 162526
rect 362542 162438 362722 162526
rect 362830 162438 363010 162526
rect 363264 162438 363444 162526
rect 363552 162438 363732 162526
rect 363840 162438 364020 162526
rect 364128 162438 364308 162526
rect 364416 162438 364596 162526
rect 364704 162438 364884 162526
rect 364992 162438 365172 162526
rect 365280 162438 365460 162526
rect 365714 162438 365894 162526
rect 366002 162438 366182 162526
rect 366290 162438 366470 162526
rect 366578 162438 366758 162526
rect 366866 162438 367046 162526
rect 367154 162438 367334 162526
rect 367442 162438 367622 162526
rect 367730 162438 367910 162526
rect 243214 162222 243394 162310
rect 243502 162222 243682 162310
rect 243790 162222 243970 162310
rect 244078 162222 244258 162310
rect 244366 162222 244546 162310
rect 244654 162222 244834 162310
rect 244942 162222 245122 162310
rect 245230 162222 245410 162310
rect 245664 162222 245844 162310
rect 245952 162222 246132 162310
rect 246240 162222 246420 162310
rect 246528 162222 246708 162310
rect 246816 162222 246996 162310
rect 247104 162222 247284 162310
rect 247392 162222 247572 162310
rect 247680 162222 247860 162310
rect 248114 162222 248294 162310
rect 248402 162222 248582 162310
rect 248690 162222 248870 162310
rect 248978 162222 249158 162310
rect 249266 162222 249446 162310
rect 249554 162222 249734 162310
rect 249842 162222 250022 162310
rect 250130 162222 250310 162310
rect 250564 162222 250744 162310
rect 360436 162222 360560 162310
rect 360814 162222 360994 162310
rect 361102 162222 361282 162310
rect 361390 162222 361570 162310
rect 361678 162222 361858 162310
rect 361966 162222 362146 162310
rect 362254 162222 362434 162310
rect 362542 162222 362722 162310
rect 362830 162222 363010 162310
rect 363264 162222 363444 162310
rect 363552 162222 363732 162310
rect 363840 162222 364020 162310
rect 364128 162222 364308 162310
rect 364416 162222 364596 162310
rect 364704 162222 364884 162310
rect 364992 162222 365172 162310
rect 365280 162222 365460 162310
rect 365714 162222 365894 162310
rect 366002 162222 366182 162310
rect 366290 162222 366470 162310
rect 366578 162222 366758 162310
rect 366866 162222 367046 162310
rect 367154 162222 367334 162310
rect 367442 162222 367622 162310
rect 367730 162222 367910 162310
rect 243214 161746 243394 161834
rect 243502 161746 243682 161834
rect 243790 161746 243970 161834
rect 244078 161746 244258 161834
rect 244366 161746 244546 161834
rect 244654 161746 244834 161834
rect 244942 161746 245122 161834
rect 245230 161746 245410 161834
rect 245664 161746 245844 161834
rect 245952 161746 246132 161834
rect 246240 161746 246420 161834
rect 246528 161746 246708 161834
rect 246816 161746 246996 161834
rect 247104 161746 247284 161834
rect 247392 161746 247572 161834
rect 247680 161746 247860 161834
rect 248114 161746 248294 161834
rect 248402 161746 248582 161834
rect 248690 161746 248870 161834
rect 248978 161746 249158 161834
rect 249266 161746 249446 161834
rect 249554 161746 249734 161834
rect 249842 161746 250022 161834
rect 250130 161746 250310 161834
rect 250564 161746 250744 161834
rect 360436 161746 360560 161834
rect 360814 161746 360994 161834
rect 361102 161746 361282 161834
rect 361390 161746 361570 161834
rect 361678 161746 361858 161834
rect 361966 161746 362146 161834
rect 362254 161746 362434 161834
rect 362542 161746 362722 161834
rect 362830 161746 363010 161834
rect 363264 161746 363444 161834
rect 363552 161746 363732 161834
rect 363840 161746 364020 161834
rect 364128 161746 364308 161834
rect 364416 161746 364596 161834
rect 364704 161746 364884 161834
rect 364992 161746 365172 161834
rect 365280 161746 365460 161834
rect 365714 161746 365894 161834
rect 366002 161746 366182 161834
rect 366290 161746 366470 161834
rect 366578 161746 366758 161834
rect 366866 161746 367046 161834
rect 367154 161746 367334 161834
rect 367442 161746 367622 161834
rect 367730 161746 367910 161834
rect 243214 161530 243394 161618
rect 243502 161530 243682 161618
rect 243790 161530 243970 161618
rect 244078 161530 244258 161618
rect 244366 161530 244546 161618
rect 244654 161530 244834 161618
rect 244942 161530 245122 161618
rect 245230 161530 245410 161618
rect 245664 161530 245844 161618
rect 245952 161530 246132 161618
rect 246240 161530 246420 161618
rect 246528 161530 246708 161618
rect 246816 161530 246996 161618
rect 247104 161530 247284 161618
rect 247392 161530 247572 161618
rect 247680 161530 247860 161618
rect 248114 161530 248294 161618
rect 248402 161530 248582 161618
rect 248690 161530 248870 161618
rect 248978 161530 249158 161618
rect 249266 161530 249446 161618
rect 249554 161530 249734 161618
rect 249842 161530 250022 161618
rect 250130 161530 250310 161618
rect 250564 161530 250744 161618
rect 360436 161530 360560 161618
rect 360814 161530 360994 161618
rect 361102 161530 361282 161618
rect 361390 161530 361570 161618
rect 361678 161530 361858 161618
rect 361966 161530 362146 161618
rect 362254 161530 362434 161618
rect 362542 161530 362722 161618
rect 362830 161530 363010 161618
rect 363264 161530 363444 161618
rect 363552 161530 363732 161618
rect 363840 161530 364020 161618
rect 364128 161530 364308 161618
rect 364416 161530 364596 161618
rect 364704 161530 364884 161618
rect 364992 161530 365172 161618
rect 365280 161530 365460 161618
rect 365714 161530 365894 161618
rect 366002 161530 366182 161618
rect 366290 161530 366470 161618
rect 366578 161530 366758 161618
rect 366866 161530 367046 161618
rect 367154 161530 367334 161618
rect 367442 161530 367622 161618
rect 367730 161530 367910 161618
rect 243214 161054 243394 161142
rect 243502 161054 243682 161142
rect 243790 161054 243970 161142
rect 244078 161054 244258 161142
rect 244366 161054 244546 161142
rect 244654 161054 244834 161142
rect 244942 161054 245122 161142
rect 245230 161054 245410 161142
rect 245664 161054 245844 161142
rect 245952 161054 246132 161142
rect 246240 161054 246420 161142
rect 246528 161054 246708 161142
rect 246816 161054 246996 161142
rect 247104 161054 247284 161142
rect 247392 161054 247572 161142
rect 247680 161054 247860 161142
rect 248114 161054 248294 161142
rect 248402 161054 248582 161142
rect 248690 161054 248870 161142
rect 248978 161054 249158 161142
rect 249266 161054 249446 161142
rect 249554 161054 249734 161142
rect 249842 161054 250022 161142
rect 250130 161054 250310 161142
rect 250564 161054 250744 161142
rect 360436 161054 360560 161142
rect 360814 161054 360994 161142
rect 361102 161054 361282 161142
rect 361390 161054 361570 161142
rect 361678 161054 361858 161142
rect 361966 161054 362146 161142
rect 362254 161054 362434 161142
rect 362542 161054 362722 161142
rect 362830 161054 363010 161142
rect 363264 161054 363444 161142
rect 363552 161054 363732 161142
rect 363840 161054 364020 161142
rect 364128 161054 364308 161142
rect 364416 161054 364596 161142
rect 364704 161054 364884 161142
rect 364992 161054 365172 161142
rect 365280 161054 365460 161142
rect 365714 161054 365894 161142
rect 366002 161054 366182 161142
rect 366290 161054 366470 161142
rect 366578 161054 366758 161142
rect 366866 161054 367046 161142
rect 367154 161054 367334 161142
rect 367442 161054 367622 161142
rect 367730 161054 367910 161142
rect 243214 160580 243394 160668
rect 243502 160580 243682 160668
rect 243790 160580 243970 160668
rect 244078 160580 244258 160668
rect 244366 160580 244546 160668
rect 244654 160580 244834 160668
rect 244942 160580 245122 160668
rect 245230 160580 245410 160668
rect 245664 160580 245844 160668
rect 245952 160580 246132 160668
rect 246240 160580 246420 160668
rect 246528 160580 246708 160668
rect 246816 160580 246996 160668
rect 247104 160580 247284 160668
rect 247392 160580 247572 160668
rect 247680 160580 247860 160668
rect 248114 160580 248294 160668
rect 248402 160580 248582 160668
rect 248690 160580 248870 160668
rect 248978 160580 249158 160668
rect 249266 160580 249446 160668
rect 249554 160580 249734 160668
rect 249842 160580 250022 160668
rect 250130 160580 250310 160668
rect 250564 160580 250744 160668
rect 360436 160580 360560 160668
rect 360814 160580 360994 160668
rect 361102 160580 361282 160668
rect 361390 160580 361570 160668
rect 361678 160580 361858 160668
rect 361966 160580 362146 160668
rect 362254 160580 362434 160668
rect 362542 160580 362722 160668
rect 362830 160580 363010 160668
rect 363264 160580 363444 160668
rect 363552 160580 363732 160668
rect 363840 160580 364020 160668
rect 364128 160580 364308 160668
rect 364416 160580 364596 160668
rect 364704 160580 364884 160668
rect 364992 160580 365172 160668
rect 365280 160580 365460 160668
rect 365714 160580 365894 160668
rect 366002 160580 366182 160668
rect 366290 160580 366470 160668
rect 366578 160580 366758 160668
rect 366866 160580 367046 160668
rect 367154 160580 367334 160668
rect 367442 160580 367622 160668
rect 367730 160580 367910 160668
rect 243214 160104 243394 160192
rect 243502 160104 243682 160192
rect 243790 160104 243970 160192
rect 244078 160104 244258 160192
rect 244366 160104 244546 160192
rect 244654 160104 244834 160192
rect 244942 160104 245122 160192
rect 245230 160104 245410 160192
rect 245664 160104 245844 160192
rect 245952 160104 246132 160192
rect 246240 160104 246420 160192
rect 246528 160104 246708 160192
rect 246816 160104 246996 160192
rect 247104 160104 247284 160192
rect 247392 160104 247572 160192
rect 247680 160104 247860 160192
rect 248114 160104 248294 160192
rect 248402 160104 248582 160192
rect 248690 160104 248870 160192
rect 248978 160104 249158 160192
rect 249266 160104 249446 160192
rect 249554 160104 249734 160192
rect 249842 160104 250022 160192
rect 250130 160104 250310 160192
rect 250564 160104 250744 160192
rect 360436 160104 360560 160192
rect 360814 160104 360994 160192
rect 361102 160104 361282 160192
rect 361390 160104 361570 160192
rect 361678 160104 361858 160192
rect 361966 160104 362146 160192
rect 362254 160104 362434 160192
rect 362542 160104 362722 160192
rect 362830 160104 363010 160192
rect 363264 160104 363444 160192
rect 363552 160104 363732 160192
rect 363840 160104 364020 160192
rect 364128 160104 364308 160192
rect 364416 160104 364596 160192
rect 364704 160104 364884 160192
rect 364992 160104 365172 160192
rect 365280 160104 365460 160192
rect 365714 160104 365894 160192
rect 366002 160104 366182 160192
rect 366290 160104 366470 160192
rect 366578 160104 366758 160192
rect 366866 160104 367046 160192
rect 367154 160104 367334 160192
rect 367442 160104 367622 160192
rect 367730 160104 367910 160192
rect 243214 159888 243394 159976
rect 243502 159888 243682 159976
rect 243790 159888 243970 159976
rect 244078 159888 244258 159976
rect 244366 159888 244546 159976
rect 244654 159888 244834 159976
rect 244942 159888 245122 159976
rect 245230 159888 245410 159976
rect 245664 159888 245844 159976
rect 245952 159888 246132 159976
rect 246240 159888 246420 159976
rect 246528 159888 246708 159976
rect 246816 159888 246996 159976
rect 247104 159888 247284 159976
rect 247392 159888 247572 159976
rect 247680 159888 247860 159976
rect 248114 159888 248294 159976
rect 248402 159888 248582 159976
rect 248690 159888 248870 159976
rect 248978 159888 249158 159976
rect 249266 159888 249446 159976
rect 249554 159888 249734 159976
rect 249842 159888 250022 159976
rect 250130 159888 250310 159976
rect 250564 159888 250744 159976
rect 360436 159888 360560 159976
rect 360814 159888 360994 159976
rect 361102 159888 361282 159976
rect 361390 159888 361570 159976
rect 361678 159888 361858 159976
rect 361966 159888 362146 159976
rect 362254 159888 362434 159976
rect 362542 159888 362722 159976
rect 362830 159888 363010 159976
rect 363264 159888 363444 159976
rect 363552 159888 363732 159976
rect 363840 159888 364020 159976
rect 364128 159888 364308 159976
rect 364416 159888 364596 159976
rect 364704 159888 364884 159976
rect 364992 159888 365172 159976
rect 365280 159888 365460 159976
rect 365714 159888 365894 159976
rect 366002 159888 366182 159976
rect 366290 159888 366470 159976
rect 366578 159888 366758 159976
rect 366866 159888 367046 159976
rect 367154 159888 367334 159976
rect 367442 159888 367622 159976
rect 367730 159888 367910 159976
rect 243214 159412 243394 159500
rect 243502 159412 243682 159500
rect 243790 159412 243970 159500
rect 244078 159412 244258 159500
rect 244366 159412 244546 159500
rect 244654 159412 244834 159500
rect 244942 159412 245122 159500
rect 245230 159412 245410 159500
rect 245664 159412 245844 159500
rect 245952 159412 246132 159500
rect 246240 159412 246420 159500
rect 246528 159412 246708 159500
rect 246816 159412 246996 159500
rect 247104 159412 247284 159500
rect 247392 159412 247572 159500
rect 247680 159412 247860 159500
rect 248114 159412 248294 159500
rect 248402 159412 248582 159500
rect 248690 159412 248870 159500
rect 248978 159412 249158 159500
rect 249266 159412 249446 159500
rect 249554 159412 249734 159500
rect 249842 159412 250022 159500
rect 250130 159412 250310 159500
rect 250564 159412 250744 159500
rect 360436 159412 360560 159500
rect 360814 159412 360994 159500
rect 361102 159412 361282 159500
rect 361390 159412 361570 159500
rect 361678 159412 361858 159500
rect 361966 159412 362146 159500
rect 362254 159412 362434 159500
rect 362542 159412 362722 159500
rect 362830 159412 363010 159500
rect 363264 159412 363444 159500
rect 363552 159412 363732 159500
rect 363840 159412 364020 159500
rect 364128 159412 364308 159500
rect 364416 159412 364596 159500
rect 364704 159412 364884 159500
rect 364992 159412 365172 159500
rect 365280 159412 365460 159500
rect 365714 159412 365894 159500
rect 366002 159412 366182 159500
rect 366290 159412 366470 159500
rect 366578 159412 366758 159500
rect 366866 159412 367046 159500
rect 367154 159412 367334 159500
rect 367442 159412 367622 159500
rect 367730 159412 367910 159500
rect 243214 159196 243394 159284
rect 243502 159196 243682 159284
rect 243790 159196 243970 159284
rect 244078 159196 244258 159284
rect 244366 159196 244546 159284
rect 244654 159196 244834 159284
rect 244942 159196 245122 159284
rect 245230 159196 245410 159284
rect 245664 159196 245844 159284
rect 245952 159196 246132 159284
rect 246240 159196 246420 159284
rect 246528 159196 246708 159284
rect 246816 159196 246996 159284
rect 247104 159196 247284 159284
rect 247392 159196 247572 159284
rect 247680 159196 247860 159284
rect 248114 159196 248294 159284
rect 248402 159196 248582 159284
rect 248690 159196 248870 159284
rect 248978 159196 249158 159284
rect 249266 159196 249446 159284
rect 249554 159196 249734 159284
rect 249842 159196 250022 159284
rect 250130 159196 250310 159284
rect 250564 159196 250744 159284
rect 360436 159196 360560 159284
rect 360814 159196 360994 159284
rect 361102 159196 361282 159284
rect 361390 159196 361570 159284
rect 361678 159196 361858 159284
rect 361966 159196 362146 159284
rect 362254 159196 362434 159284
rect 362542 159196 362722 159284
rect 362830 159196 363010 159284
rect 363264 159196 363444 159284
rect 363552 159196 363732 159284
rect 363840 159196 364020 159284
rect 364128 159196 364308 159284
rect 364416 159196 364596 159284
rect 364704 159196 364884 159284
rect 364992 159196 365172 159284
rect 365280 159196 365460 159284
rect 365714 159196 365894 159284
rect 366002 159196 366182 159284
rect 366290 159196 366470 159284
rect 366578 159196 366758 159284
rect 366866 159196 367046 159284
rect 367154 159196 367334 159284
rect 367442 159196 367622 159284
rect 367730 159196 367910 159284
rect 243214 158720 243394 158808
rect 243502 158720 243682 158808
rect 243790 158720 243970 158808
rect 244078 158720 244258 158808
rect 244366 158720 244546 158808
rect 244654 158720 244834 158808
rect 244942 158720 245122 158808
rect 245230 158720 245410 158808
rect 245664 158720 245844 158808
rect 245952 158720 246132 158808
rect 246240 158720 246420 158808
rect 246528 158720 246708 158808
rect 246816 158720 246996 158808
rect 247104 158720 247284 158808
rect 247392 158720 247572 158808
rect 247680 158720 247860 158808
rect 248114 158720 248294 158808
rect 248402 158720 248582 158808
rect 248690 158720 248870 158808
rect 248978 158720 249158 158808
rect 249266 158720 249446 158808
rect 249554 158720 249734 158808
rect 249842 158720 250022 158808
rect 250130 158720 250310 158808
rect 250564 158720 250744 158808
rect 360436 158720 360560 158808
rect 360814 158720 360994 158808
rect 361102 158720 361282 158808
rect 361390 158720 361570 158808
rect 361678 158720 361858 158808
rect 361966 158720 362146 158808
rect 362254 158720 362434 158808
rect 362542 158720 362722 158808
rect 362830 158720 363010 158808
rect 363264 158720 363444 158808
rect 363552 158720 363732 158808
rect 363840 158720 364020 158808
rect 364128 158720 364308 158808
rect 364416 158720 364596 158808
rect 364704 158720 364884 158808
rect 364992 158720 365172 158808
rect 365280 158720 365460 158808
rect 365714 158720 365894 158808
rect 366002 158720 366182 158808
rect 366290 158720 366470 158808
rect 366578 158720 366758 158808
rect 366866 158720 367046 158808
rect 367154 158720 367334 158808
rect 367442 158720 367622 158808
rect 367730 158720 367910 158808
rect 243214 158504 243394 158592
rect 243502 158504 243682 158592
rect 243790 158504 243970 158592
rect 244078 158504 244258 158592
rect 244366 158504 244546 158592
rect 244654 158504 244834 158592
rect 244942 158504 245122 158592
rect 245230 158504 245410 158592
rect 245664 158504 245844 158592
rect 245952 158504 246132 158592
rect 246240 158504 246420 158592
rect 246528 158504 246708 158592
rect 246816 158504 246996 158592
rect 247104 158504 247284 158592
rect 247392 158504 247572 158592
rect 247680 158504 247860 158592
rect 248114 158504 248294 158592
rect 248402 158504 248582 158592
rect 248690 158504 248870 158592
rect 248978 158504 249158 158592
rect 249266 158504 249446 158592
rect 249554 158504 249734 158592
rect 249842 158504 250022 158592
rect 250130 158504 250310 158592
rect 250564 158504 250744 158592
rect 360436 158504 360560 158592
rect 360814 158504 360994 158592
rect 361102 158504 361282 158592
rect 361390 158504 361570 158592
rect 361678 158504 361858 158592
rect 361966 158504 362146 158592
rect 362254 158504 362434 158592
rect 362542 158504 362722 158592
rect 362830 158504 363010 158592
rect 363264 158504 363444 158592
rect 363552 158504 363732 158592
rect 363840 158504 364020 158592
rect 364128 158504 364308 158592
rect 364416 158504 364596 158592
rect 364704 158504 364884 158592
rect 364992 158504 365172 158592
rect 365280 158504 365460 158592
rect 365714 158504 365894 158592
rect 366002 158504 366182 158592
rect 366290 158504 366470 158592
rect 366578 158504 366758 158592
rect 366866 158504 367046 158592
rect 367154 158504 367334 158592
rect 367442 158504 367622 158592
rect 367730 158504 367910 158592
rect 243214 158028 243394 158116
rect 243502 158028 243682 158116
rect 243790 158028 243970 158116
rect 244078 158028 244258 158116
rect 244366 158028 244546 158116
rect 244654 158028 244834 158116
rect 244942 158028 245122 158116
rect 245230 158028 245410 158116
rect 245664 158028 245844 158116
rect 245952 158028 246132 158116
rect 246240 158028 246420 158116
rect 246528 158028 246708 158116
rect 246816 158028 246996 158116
rect 247104 158028 247284 158116
rect 247392 158028 247572 158116
rect 247680 158028 247860 158116
rect 248114 158028 248294 158116
rect 248402 158028 248582 158116
rect 248690 158028 248870 158116
rect 248978 158028 249158 158116
rect 249266 158028 249446 158116
rect 249554 158028 249734 158116
rect 249842 158028 250022 158116
rect 250130 158028 250310 158116
rect 250564 158028 250744 158116
rect 360436 158028 360560 158116
rect 360814 158028 360994 158116
rect 361102 158028 361282 158116
rect 361390 158028 361570 158116
rect 361678 158028 361858 158116
rect 361966 158028 362146 158116
rect 362254 158028 362434 158116
rect 362542 158028 362722 158116
rect 362830 158028 363010 158116
rect 363264 158028 363444 158116
rect 363552 158028 363732 158116
rect 363840 158028 364020 158116
rect 364128 158028 364308 158116
rect 364416 158028 364596 158116
rect 364704 158028 364884 158116
rect 364992 158028 365172 158116
rect 365280 158028 365460 158116
rect 365714 158028 365894 158116
rect 366002 158028 366182 158116
rect 366290 158028 366470 158116
rect 366578 158028 366758 158116
rect 366866 158028 367046 158116
rect 367154 158028 367334 158116
rect 367442 158028 367622 158116
rect 367730 158028 367910 158116
rect 243214 157554 243394 157642
rect 243502 157554 243682 157642
rect 243790 157554 243970 157642
rect 244078 157554 244258 157642
rect 244366 157554 244546 157642
rect 244654 157554 244834 157642
rect 244942 157554 245122 157642
rect 245230 157554 245410 157642
rect 245664 157554 245844 157642
rect 245952 157554 246132 157642
rect 246240 157554 246420 157642
rect 246528 157554 246708 157642
rect 246816 157554 246996 157642
rect 247104 157554 247284 157642
rect 247392 157554 247572 157642
rect 247680 157554 247860 157642
rect 248114 157554 248294 157642
rect 248402 157554 248582 157642
rect 248690 157554 248870 157642
rect 248978 157554 249158 157642
rect 249266 157554 249446 157642
rect 249554 157554 249734 157642
rect 249842 157554 250022 157642
rect 250130 157554 250310 157642
rect 250564 157554 250744 157642
rect 360436 157554 360560 157642
rect 360814 157554 360994 157642
rect 361102 157554 361282 157642
rect 361390 157554 361570 157642
rect 361678 157554 361858 157642
rect 361966 157554 362146 157642
rect 362254 157554 362434 157642
rect 362542 157554 362722 157642
rect 362830 157554 363010 157642
rect 363264 157554 363444 157642
rect 363552 157554 363732 157642
rect 363840 157554 364020 157642
rect 364128 157554 364308 157642
rect 364416 157554 364596 157642
rect 364704 157554 364884 157642
rect 364992 157554 365172 157642
rect 365280 157554 365460 157642
rect 365714 157554 365894 157642
rect 366002 157554 366182 157642
rect 366290 157554 366470 157642
rect 366578 157554 366758 157642
rect 366866 157554 367046 157642
rect 367154 157554 367334 157642
rect 367442 157554 367622 157642
rect 367730 157554 367910 157642
rect 243214 157078 243394 157166
rect 243502 157078 243682 157166
rect 243790 157078 243970 157166
rect 244078 157078 244258 157166
rect 244366 157078 244546 157166
rect 244654 157078 244834 157166
rect 244942 157078 245122 157166
rect 245230 157078 245410 157166
rect 245664 157078 245844 157166
rect 245952 157078 246132 157166
rect 246240 157078 246420 157166
rect 246528 157078 246708 157166
rect 246816 157078 246996 157166
rect 247104 157078 247284 157166
rect 247392 157078 247572 157166
rect 247680 157078 247860 157166
rect 248114 157078 248294 157166
rect 248402 157078 248582 157166
rect 248690 157078 248870 157166
rect 248978 157078 249158 157166
rect 249266 157078 249446 157166
rect 249554 157078 249734 157166
rect 249842 157078 250022 157166
rect 250130 157078 250310 157166
rect 250564 157078 250744 157166
rect 360436 157078 360560 157166
rect 360814 157078 360994 157166
rect 361102 157078 361282 157166
rect 361390 157078 361570 157166
rect 361678 157078 361858 157166
rect 361966 157078 362146 157166
rect 362254 157078 362434 157166
rect 362542 157078 362722 157166
rect 362830 157078 363010 157166
rect 363264 157078 363444 157166
rect 363552 157078 363732 157166
rect 363840 157078 364020 157166
rect 364128 157078 364308 157166
rect 364416 157078 364596 157166
rect 364704 157078 364884 157166
rect 364992 157078 365172 157166
rect 365280 157078 365460 157166
rect 365714 157078 365894 157166
rect 366002 157078 366182 157166
rect 366290 157078 366470 157166
rect 366578 157078 366758 157166
rect 366866 157078 367046 157166
rect 367154 157078 367334 157166
rect 367442 157078 367622 157166
rect 367730 157078 367910 157166
rect 243214 156862 243394 156950
rect 243502 156862 243682 156950
rect 243790 156862 243970 156950
rect 244078 156862 244258 156950
rect 244366 156862 244546 156950
rect 244654 156862 244834 156950
rect 244942 156862 245122 156950
rect 245230 156862 245410 156950
rect 245664 156862 245844 156950
rect 245952 156862 246132 156950
rect 246240 156862 246420 156950
rect 246528 156862 246708 156950
rect 246816 156862 246996 156950
rect 247104 156862 247284 156950
rect 247392 156862 247572 156950
rect 247680 156862 247860 156950
rect 248114 156862 248294 156950
rect 248402 156862 248582 156950
rect 248690 156862 248870 156950
rect 248978 156862 249158 156950
rect 249266 156862 249446 156950
rect 249554 156862 249734 156950
rect 249842 156862 250022 156950
rect 250130 156862 250310 156950
rect 250564 156862 250744 156950
rect 360436 156862 360560 156950
rect 360814 156862 360994 156950
rect 361102 156862 361282 156950
rect 361390 156862 361570 156950
rect 361678 156862 361858 156950
rect 361966 156862 362146 156950
rect 362254 156862 362434 156950
rect 362542 156862 362722 156950
rect 362830 156862 363010 156950
rect 363264 156862 363444 156950
rect 363552 156862 363732 156950
rect 363840 156862 364020 156950
rect 364128 156862 364308 156950
rect 364416 156862 364596 156950
rect 364704 156862 364884 156950
rect 364992 156862 365172 156950
rect 365280 156862 365460 156950
rect 365714 156862 365894 156950
rect 366002 156862 366182 156950
rect 366290 156862 366470 156950
rect 366578 156862 366758 156950
rect 366866 156862 367046 156950
rect 367154 156862 367334 156950
rect 367442 156862 367622 156950
rect 367730 156862 367910 156950
rect 243214 156386 243394 156474
rect 243502 156386 243682 156474
rect 243790 156386 243970 156474
rect 244078 156386 244258 156474
rect 244366 156386 244546 156474
rect 244654 156386 244834 156474
rect 244942 156386 245122 156474
rect 245230 156386 245410 156474
rect 245664 156386 245844 156474
rect 245952 156386 246132 156474
rect 246240 156386 246420 156474
rect 246528 156386 246708 156474
rect 246816 156386 246996 156474
rect 247104 156386 247284 156474
rect 247392 156386 247572 156474
rect 247680 156386 247860 156474
rect 248114 156386 248294 156474
rect 248402 156386 248582 156474
rect 248690 156386 248870 156474
rect 248978 156386 249158 156474
rect 249266 156386 249446 156474
rect 249554 156386 249734 156474
rect 249842 156386 250022 156474
rect 250130 156386 250310 156474
rect 250564 156386 250744 156474
rect 360436 156386 360560 156474
rect 360814 156386 360994 156474
rect 361102 156386 361282 156474
rect 361390 156386 361570 156474
rect 361678 156386 361858 156474
rect 361966 156386 362146 156474
rect 362254 156386 362434 156474
rect 362542 156386 362722 156474
rect 362830 156386 363010 156474
rect 363264 156386 363444 156474
rect 363552 156386 363732 156474
rect 363840 156386 364020 156474
rect 364128 156386 364308 156474
rect 364416 156386 364596 156474
rect 364704 156386 364884 156474
rect 364992 156386 365172 156474
rect 365280 156386 365460 156474
rect 365714 156386 365894 156474
rect 366002 156386 366182 156474
rect 366290 156386 366470 156474
rect 366578 156386 366758 156474
rect 366866 156386 367046 156474
rect 367154 156386 367334 156474
rect 367442 156386 367622 156474
rect 367730 156386 367910 156474
rect 243214 156170 243394 156258
rect 243502 156170 243682 156258
rect 243790 156170 243970 156258
rect 244078 156170 244258 156258
rect 244366 156170 244546 156258
rect 244654 156170 244834 156258
rect 244942 156170 245122 156258
rect 245230 156170 245410 156258
rect 245664 156170 245844 156258
rect 245952 156170 246132 156258
rect 246240 156170 246420 156258
rect 246528 156170 246708 156258
rect 246816 156170 246996 156258
rect 247104 156170 247284 156258
rect 247392 156170 247572 156258
rect 247680 156170 247860 156258
rect 248114 156170 248294 156258
rect 248402 156170 248582 156258
rect 248690 156170 248870 156258
rect 248978 156170 249158 156258
rect 249266 156170 249446 156258
rect 249554 156170 249734 156258
rect 249842 156170 250022 156258
rect 250130 156170 250310 156258
rect 250564 156170 250744 156258
rect 360436 156170 360560 156258
rect 360814 156170 360994 156258
rect 361102 156170 361282 156258
rect 361390 156170 361570 156258
rect 361678 156170 361858 156258
rect 361966 156170 362146 156258
rect 362254 156170 362434 156258
rect 362542 156170 362722 156258
rect 362830 156170 363010 156258
rect 363264 156170 363444 156258
rect 363552 156170 363732 156258
rect 363840 156170 364020 156258
rect 364128 156170 364308 156258
rect 364416 156170 364596 156258
rect 364704 156170 364884 156258
rect 364992 156170 365172 156258
rect 365280 156170 365460 156258
rect 365714 156170 365894 156258
rect 366002 156170 366182 156258
rect 366290 156170 366470 156258
rect 366578 156170 366758 156258
rect 366866 156170 367046 156258
rect 367154 156170 367334 156258
rect 367442 156170 367622 156258
rect 367730 156170 367910 156258
rect 243214 155694 243394 155782
rect 243502 155694 243682 155782
rect 243790 155694 243970 155782
rect 244078 155694 244258 155782
rect 244366 155694 244546 155782
rect 244654 155694 244834 155782
rect 244942 155694 245122 155782
rect 245230 155694 245410 155782
rect 245664 155694 245844 155782
rect 245952 155694 246132 155782
rect 246240 155694 246420 155782
rect 246528 155694 246708 155782
rect 246816 155694 246996 155782
rect 247104 155694 247284 155782
rect 247392 155694 247572 155782
rect 247680 155694 247860 155782
rect 248114 155694 248294 155782
rect 248402 155694 248582 155782
rect 248690 155694 248870 155782
rect 248978 155694 249158 155782
rect 249266 155694 249446 155782
rect 249554 155694 249734 155782
rect 249842 155694 250022 155782
rect 250130 155694 250310 155782
rect 250564 155694 250744 155782
rect 360436 155694 360560 155782
rect 360814 155694 360994 155782
rect 361102 155694 361282 155782
rect 361390 155694 361570 155782
rect 361678 155694 361858 155782
rect 361966 155694 362146 155782
rect 362254 155694 362434 155782
rect 362542 155694 362722 155782
rect 362830 155694 363010 155782
rect 363264 155694 363444 155782
rect 363552 155694 363732 155782
rect 363840 155694 364020 155782
rect 364128 155694 364308 155782
rect 364416 155694 364596 155782
rect 364704 155694 364884 155782
rect 364992 155694 365172 155782
rect 365280 155694 365460 155782
rect 365714 155694 365894 155782
rect 366002 155694 366182 155782
rect 366290 155694 366470 155782
rect 366578 155694 366758 155782
rect 366866 155694 367046 155782
rect 367154 155694 367334 155782
rect 367442 155694 367622 155782
rect 367730 155694 367910 155782
rect 243214 155478 243394 155566
rect 243502 155478 243682 155566
rect 243790 155478 243970 155566
rect 244078 155478 244258 155566
rect 244366 155478 244546 155566
rect 244654 155478 244834 155566
rect 244942 155478 245122 155566
rect 245230 155478 245410 155566
rect 245664 155478 245844 155566
rect 245952 155478 246132 155566
rect 246240 155478 246420 155566
rect 246528 155478 246708 155566
rect 246816 155478 246996 155566
rect 247104 155478 247284 155566
rect 247392 155478 247572 155566
rect 247680 155478 247860 155566
rect 248114 155478 248294 155566
rect 248402 155478 248582 155566
rect 248690 155478 248870 155566
rect 248978 155478 249158 155566
rect 249266 155478 249446 155566
rect 249554 155478 249734 155566
rect 249842 155478 250022 155566
rect 250130 155478 250310 155566
rect 250564 155478 250744 155566
rect 360436 155478 360560 155566
rect 360814 155478 360994 155566
rect 361102 155478 361282 155566
rect 361390 155478 361570 155566
rect 361678 155478 361858 155566
rect 361966 155478 362146 155566
rect 362254 155478 362434 155566
rect 362542 155478 362722 155566
rect 362830 155478 363010 155566
rect 363264 155478 363444 155566
rect 363552 155478 363732 155566
rect 363840 155478 364020 155566
rect 364128 155478 364308 155566
rect 364416 155478 364596 155566
rect 364704 155478 364884 155566
rect 364992 155478 365172 155566
rect 365280 155478 365460 155566
rect 365714 155478 365894 155566
rect 366002 155478 366182 155566
rect 366290 155478 366470 155566
rect 366578 155478 366758 155566
rect 366866 155478 367046 155566
rect 367154 155478 367334 155566
rect 367442 155478 367622 155566
rect 367730 155478 367910 155566
rect 243214 155002 243394 155090
rect 243502 155002 243682 155090
rect 243790 155002 243970 155090
rect 244078 155002 244258 155090
rect 244366 155002 244546 155090
rect 244654 155002 244834 155090
rect 244942 155002 245122 155090
rect 245230 155002 245410 155090
rect 245664 155002 245844 155090
rect 245952 155002 246132 155090
rect 246240 155002 246420 155090
rect 246528 155002 246708 155090
rect 246816 155002 246996 155090
rect 247104 155002 247284 155090
rect 247392 155002 247572 155090
rect 247680 155002 247860 155090
rect 248114 155002 248294 155090
rect 248402 155002 248582 155090
rect 248690 155002 248870 155090
rect 248978 155002 249158 155090
rect 249266 155002 249446 155090
rect 249554 155002 249734 155090
rect 249842 155002 250022 155090
rect 250130 155002 250310 155090
rect 250564 155002 250744 155090
rect 360436 155002 360560 155090
rect 360814 155002 360994 155090
rect 361102 155002 361282 155090
rect 361390 155002 361570 155090
rect 361678 155002 361858 155090
rect 361966 155002 362146 155090
rect 362254 155002 362434 155090
rect 362542 155002 362722 155090
rect 362830 155002 363010 155090
rect 363264 155002 363444 155090
rect 363552 155002 363732 155090
rect 363840 155002 364020 155090
rect 364128 155002 364308 155090
rect 364416 155002 364596 155090
rect 364704 155002 364884 155090
rect 364992 155002 365172 155090
rect 365280 155002 365460 155090
rect 365714 155002 365894 155090
rect 366002 155002 366182 155090
rect 366290 155002 366470 155090
rect 366578 155002 366758 155090
rect 366866 155002 367046 155090
rect 367154 155002 367334 155090
rect 367442 155002 367622 155090
rect 367730 155002 367910 155090
rect 243214 154528 243394 154616
rect 243502 154528 243682 154616
rect 243790 154528 243970 154616
rect 244078 154528 244258 154616
rect 244366 154528 244546 154616
rect 244654 154528 244834 154616
rect 244942 154528 245122 154616
rect 245230 154528 245410 154616
rect 245664 154528 245844 154616
rect 245952 154528 246132 154616
rect 246240 154528 246420 154616
rect 246528 154528 246708 154616
rect 246816 154528 246996 154616
rect 247104 154528 247284 154616
rect 247392 154528 247572 154616
rect 247680 154528 247860 154616
rect 248114 154528 248294 154616
rect 248402 154528 248582 154616
rect 248690 154528 248870 154616
rect 248978 154528 249158 154616
rect 249266 154528 249446 154616
rect 249554 154528 249734 154616
rect 249842 154528 250022 154616
rect 250130 154528 250310 154616
rect 250564 154528 250744 154616
rect 360436 154528 360560 154616
rect 360814 154528 360994 154616
rect 361102 154528 361282 154616
rect 361390 154528 361570 154616
rect 361678 154528 361858 154616
rect 361966 154528 362146 154616
rect 362254 154528 362434 154616
rect 362542 154528 362722 154616
rect 362830 154528 363010 154616
rect 363264 154528 363444 154616
rect 363552 154528 363732 154616
rect 363840 154528 364020 154616
rect 364128 154528 364308 154616
rect 364416 154528 364596 154616
rect 364704 154528 364884 154616
rect 364992 154528 365172 154616
rect 365280 154528 365460 154616
rect 365714 154528 365894 154616
rect 366002 154528 366182 154616
rect 366290 154528 366470 154616
rect 366578 154528 366758 154616
rect 366866 154528 367046 154616
rect 367154 154528 367334 154616
rect 367442 154528 367622 154616
rect 367730 154528 367910 154616
rect 243214 154052 243394 154140
rect 243502 154052 243682 154140
rect 243790 154052 243970 154140
rect 244078 154052 244258 154140
rect 244366 154052 244546 154140
rect 244654 154052 244834 154140
rect 244942 154052 245122 154140
rect 245230 154052 245410 154140
rect 245664 154052 245844 154140
rect 245952 154052 246132 154140
rect 246240 154052 246420 154140
rect 246528 154052 246708 154140
rect 246816 154052 246996 154140
rect 247104 154052 247284 154140
rect 247392 154052 247572 154140
rect 247680 154052 247860 154140
rect 248114 154052 248294 154140
rect 248402 154052 248582 154140
rect 248690 154052 248870 154140
rect 248978 154052 249158 154140
rect 249266 154052 249446 154140
rect 249554 154052 249734 154140
rect 249842 154052 250022 154140
rect 250130 154052 250310 154140
rect 250564 154052 250744 154140
rect 360436 154052 360560 154140
rect 360814 154052 360994 154140
rect 361102 154052 361282 154140
rect 361390 154052 361570 154140
rect 361678 154052 361858 154140
rect 361966 154052 362146 154140
rect 362254 154052 362434 154140
rect 362542 154052 362722 154140
rect 362830 154052 363010 154140
rect 363264 154052 363444 154140
rect 363552 154052 363732 154140
rect 363840 154052 364020 154140
rect 364128 154052 364308 154140
rect 364416 154052 364596 154140
rect 364704 154052 364884 154140
rect 364992 154052 365172 154140
rect 365280 154052 365460 154140
rect 365714 154052 365894 154140
rect 366002 154052 366182 154140
rect 366290 154052 366470 154140
rect 366578 154052 366758 154140
rect 366866 154052 367046 154140
rect 367154 154052 367334 154140
rect 367442 154052 367622 154140
rect 367730 154052 367910 154140
rect 243214 153836 243394 153924
rect 243502 153836 243682 153924
rect 243790 153836 243970 153924
rect 244078 153836 244258 153924
rect 244366 153836 244546 153924
rect 244654 153836 244834 153924
rect 244942 153836 245122 153924
rect 245230 153836 245410 153924
rect 245664 153836 245844 153924
rect 245952 153836 246132 153924
rect 246240 153836 246420 153924
rect 246528 153836 246708 153924
rect 246816 153836 246996 153924
rect 247104 153836 247284 153924
rect 247392 153836 247572 153924
rect 247680 153836 247860 153924
rect 248114 153836 248294 153924
rect 248402 153836 248582 153924
rect 248690 153836 248870 153924
rect 248978 153836 249158 153924
rect 249266 153836 249446 153924
rect 249554 153836 249734 153924
rect 249842 153836 250022 153924
rect 250130 153836 250310 153924
rect 250564 153836 250744 153924
rect 360436 153836 360560 153924
rect 360814 153836 360994 153924
rect 361102 153836 361282 153924
rect 361390 153836 361570 153924
rect 361678 153836 361858 153924
rect 361966 153836 362146 153924
rect 362254 153836 362434 153924
rect 362542 153836 362722 153924
rect 362830 153836 363010 153924
rect 363264 153836 363444 153924
rect 363552 153836 363732 153924
rect 363840 153836 364020 153924
rect 364128 153836 364308 153924
rect 364416 153836 364596 153924
rect 364704 153836 364884 153924
rect 364992 153836 365172 153924
rect 365280 153836 365460 153924
rect 365714 153836 365894 153924
rect 366002 153836 366182 153924
rect 366290 153836 366470 153924
rect 366578 153836 366758 153924
rect 366866 153836 367046 153924
rect 367154 153836 367334 153924
rect 367442 153836 367622 153924
rect 367730 153836 367910 153924
rect 243214 153360 243394 153448
rect 243502 153360 243682 153448
rect 243790 153360 243970 153448
rect 244078 153360 244258 153448
rect 244366 153360 244546 153448
rect 244654 153360 244834 153448
rect 244942 153360 245122 153448
rect 245230 153360 245410 153448
rect 245664 153360 245844 153448
rect 245952 153360 246132 153448
rect 246240 153360 246420 153448
rect 246528 153360 246708 153448
rect 246816 153360 246996 153448
rect 247104 153360 247284 153448
rect 247392 153360 247572 153448
rect 247680 153360 247860 153448
rect 248114 153360 248294 153448
rect 248402 153360 248582 153448
rect 248690 153360 248870 153448
rect 248978 153360 249158 153448
rect 249266 153360 249446 153448
rect 249554 153360 249734 153448
rect 249842 153360 250022 153448
rect 250130 153360 250310 153448
rect 250564 153360 250744 153448
rect 360436 153360 360560 153448
rect 360814 153360 360994 153448
rect 361102 153360 361282 153448
rect 361390 153360 361570 153448
rect 361678 153360 361858 153448
rect 361966 153360 362146 153448
rect 362254 153360 362434 153448
rect 362542 153360 362722 153448
rect 362830 153360 363010 153448
rect 363264 153360 363444 153448
rect 363552 153360 363732 153448
rect 363840 153360 364020 153448
rect 364128 153360 364308 153448
rect 364416 153360 364596 153448
rect 364704 153360 364884 153448
rect 364992 153360 365172 153448
rect 365280 153360 365460 153448
rect 365714 153360 365894 153448
rect 366002 153360 366182 153448
rect 366290 153360 366470 153448
rect 366578 153360 366758 153448
rect 366866 153360 367046 153448
rect 367154 153360 367334 153448
rect 367442 153360 367622 153448
rect 367730 153360 367910 153448
rect 243214 153144 243394 153232
rect 243502 153144 243682 153232
rect 243790 153144 243970 153232
rect 244078 153144 244258 153232
rect 244366 153144 244546 153232
rect 244654 153144 244834 153232
rect 244942 153144 245122 153232
rect 245230 153144 245410 153232
rect 245664 153144 245844 153232
rect 245952 153144 246132 153232
rect 246240 153144 246420 153232
rect 246528 153144 246708 153232
rect 246816 153144 246996 153232
rect 247104 153144 247284 153232
rect 247392 153144 247572 153232
rect 247680 153144 247860 153232
rect 248114 153144 248294 153232
rect 248402 153144 248582 153232
rect 248690 153144 248870 153232
rect 248978 153144 249158 153232
rect 249266 153144 249446 153232
rect 249554 153144 249734 153232
rect 249842 153144 250022 153232
rect 250130 153144 250310 153232
rect 250564 153144 250744 153232
rect 360436 153144 360560 153232
rect 360814 153144 360994 153232
rect 361102 153144 361282 153232
rect 361390 153144 361570 153232
rect 361678 153144 361858 153232
rect 361966 153144 362146 153232
rect 362254 153144 362434 153232
rect 362542 153144 362722 153232
rect 362830 153144 363010 153232
rect 363264 153144 363444 153232
rect 363552 153144 363732 153232
rect 363840 153144 364020 153232
rect 364128 153144 364308 153232
rect 364416 153144 364596 153232
rect 364704 153144 364884 153232
rect 364992 153144 365172 153232
rect 365280 153144 365460 153232
rect 365714 153144 365894 153232
rect 366002 153144 366182 153232
rect 366290 153144 366470 153232
rect 366578 153144 366758 153232
rect 366866 153144 367046 153232
rect 367154 153144 367334 153232
rect 367442 153144 367622 153232
rect 367730 153144 367910 153232
rect 243214 152668 243394 152756
rect 243502 152668 243682 152756
rect 243790 152668 243970 152756
rect 244078 152668 244258 152756
rect 244366 152668 244546 152756
rect 244654 152668 244834 152756
rect 244942 152668 245122 152756
rect 245230 152668 245410 152756
rect 245664 152668 245844 152756
rect 245952 152668 246132 152756
rect 246240 152668 246420 152756
rect 246528 152668 246708 152756
rect 246816 152668 246996 152756
rect 247104 152668 247284 152756
rect 247392 152668 247572 152756
rect 247680 152668 247860 152756
rect 248114 152668 248294 152756
rect 248402 152668 248582 152756
rect 248690 152668 248870 152756
rect 248978 152668 249158 152756
rect 249266 152668 249446 152756
rect 249554 152668 249734 152756
rect 249842 152668 250022 152756
rect 250130 152668 250310 152756
rect 250564 152668 250744 152756
rect 360436 152668 360560 152756
rect 360814 152668 360994 152756
rect 361102 152668 361282 152756
rect 361390 152668 361570 152756
rect 361678 152668 361858 152756
rect 361966 152668 362146 152756
rect 362254 152668 362434 152756
rect 362542 152668 362722 152756
rect 362830 152668 363010 152756
rect 363264 152668 363444 152756
rect 363552 152668 363732 152756
rect 363840 152668 364020 152756
rect 364128 152668 364308 152756
rect 364416 152668 364596 152756
rect 364704 152668 364884 152756
rect 364992 152668 365172 152756
rect 365280 152668 365460 152756
rect 365714 152668 365894 152756
rect 366002 152668 366182 152756
rect 366290 152668 366470 152756
rect 366578 152668 366758 152756
rect 366866 152668 367046 152756
rect 367154 152668 367334 152756
rect 367442 152668 367622 152756
rect 367730 152668 367910 152756
rect 243214 152452 243394 152540
rect 243502 152452 243682 152540
rect 243790 152452 243970 152540
rect 244078 152452 244258 152540
rect 244366 152452 244546 152540
rect 244654 152452 244834 152540
rect 244942 152452 245122 152540
rect 245230 152452 245410 152540
rect 245664 152452 245844 152540
rect 245952 152452 246132 152540
rect 246240 152452 246420 152540
rect 246528 152452 246708 152540
rect 246816 152452 246996 152540
rect 247104 152452 247284 152540
rect 247392 152452 247572 152540
rect 247680 152452 247860 152540
rect 248114 152452 248294 152540
rect 248402 152452 248582 152540
rect 248690 152452 248870 152540
rect 248978 152452 249158 152540
rect 249266 152452 249446 152540
rect 249554 152452 249734 152540
rect 249842 152452 250022 152540
rect 250130 152452 250310 152540
rect 250564 152452 250744 152540
rect 360436 152452 360560 152540
rect 360814 152452 360994 152540
rect 361102 152452 361282 152540
rect 361390 152452 361570 152540
rect 361678 152452 361858 152540
rect 361966 152452 362146 152540
rect 362254 152452 362434 152540
rect 362542 152452 362722 152540
rect 362830 152452 363010 152540
rect 363264 152452 363444 152540
rect 363552 152452 363732 152540
rect 363840 152452 364020 152540
rect 364128 152452 364308 152540
rect 364416 152452 364596 152540
rect 364704 152452 364884 152540
rect 364992 152452 365172 152540
rect 365280 152452 365460 152540
rect 365714 152452 365894 152540
rect 366002 152452 366182 152540
rect 366290 152452 366470 152540
rect 366578 152452 366758 152540
rect 366866 152452 367046 152540
rect 367154 152452 367334 152540
rect 367442 152452 367622 152540
rect 367730 152452 367910 152540
rect 243214 151976 243394 152064
rect 243502 151976 243682 152064
rect 243790 151976 243970 152064
rect 244078 151976 244258 152064
rect 244366 151976 244546 152064
rect 244654 151976 244834 152064
rect 244942 151976 245122 152064
rect 245230 151976 245410 152064
rect 245664 151976 245844 152064
rect 245952 151976 246132 152064
rect 246240 151976 246420 152064
rect 246528 151976 246708 152064
rect 246816 151976 246996 152064
rect 247104 151976 247284 152064
rect 247392 151976 247572 152064
rect 247680 151976 247860 152064
rect 248114 151976 248294 152064
rect 248402 151976 248582 152064
rect 248690 151976 248870 152064
rect 248978 151976 249158 152064
rect 249266 151976 249446 152064
rect 249554 151976 249734 152064
rect 249842 151976 250022 152064
rect 250130 151976 250310 152064
rect 250564 151976 250744 152064
rect 360436 151976 360560 152064
rect 360814 151976 360994 152064
rect 361102 151976 361282 152064
rect 361390 151976 361570 152064
rect 361678 151976 361858 152064
rect 361966 151976 362146 152064
rect 362254 151976 362434 152064
rect 362542 151976 362722 152064
rect 362830 151976 363010 152064
rect 363264 151976 363444 152064
rect 363552 151976 363732 152064
rect 363840 151976 364020 152064
rect 364128 151976 364308 152064
rect 364416 151976 364596 152064
rect 364704 151976 364884 152064
rect 364992 151976 365172 152064
rect 365280 151976 365460 152064
rect 365714 151976 365894 152064
rect 366002 151976 366182 152064
rect 366290 151976 366470 152064
rect 366578 151976 366758 152064
rect 366866 151976 367046 152064
rect 367154 151976 367334 152064
rect 367442 151976 367622 152064
rect 367730 151976 367910 152064
rect 243214 151502 243394 151590
rect 243502 151502 243682 151590
rect 243790 151502 243970 151590
rect 244078 151502 244258 151590
rect 244366 151502 244546 151590
rect 244654 151502 244834 151590
rect 244942 151502 245122 151590
rect 245230 151502 245410 151590
rect 245664 151502 245844 151590
rect 245952 151502 246132 151590
rect 246240 151502 246420 151590
rect 246528 151502 246708 151590
rect 246816 151502 246996 151590
rect 247104 151502 247284 151590
rect 247392 151502 247572 151590
rect 247680 151502 247860 151590
rect 248114 151502 248294 151590
rect 248402 151502 248582 151590
rect 248690 151502 248870 151590
rect 248978 151502 249158 151590
rect 249266 151502 249446 151590
rect 249554 151502 249734 151590
rect 249842 151502 250022 151590
rect 250130 151502 250310 151590
rect 250564 151502 250744 151590
rect 360436 151502 360560 151590
rect 360814 151502 360994 151590
rect 361102 151502 361282 151590
rect 361390 151502 361570 151590
rect 361678 151502 361858 151590
rect 361966 151502 362146 151590
rect 362254 151502 362434 151590
rect 362542 151502 362722 151590
rect 362830 151502 363010 151590
rect 363264 151502 363444 151590
rect 363552 151502 363732 151590
rect 363840 151502 364020 151590
rect 364128 151502 364308 151590
rect 364416 151502 364596 151590
rect 364704 151502 364884 151590
rect 364992 151502 365172 151590
rect 365280 151502 365460 151590
rect 365714 151502 365894 151590
rect 366002 151502 366182 151590
rect 366290 151502 366470 151590
rect 366578 151502 366758 151590
rect 366866 151502 367046 151590
rect 367154 151502 367334 151590
rect 367442 151502 367622 151590
rect 367730 151502 367910 151590
rect 243214 151026 243394 151114
rect 243502 151026 243682 151114
rect 243790 151026 243970 151114
rect 244078 151026 244258 151114
rect 244366 151026 244546 151114
rect 244654 151026 244834 151114
rect 244942 151026 245122 151114
rect 245230 151026 245410 151114
rect 245664 151026 245844 151114
rect 245952 151026 246132 151114
rect 246240 151026 246420 151114
rect 246528 151026 246708 151114
rect 246816 151026 246996 151114
rect 247104 151026 247284 151114
rect 247392 151026 247572 151114
rect 247680 151026 247860 151114
rect 248114 151026 248294 151114
rect 248402 151026 248582 151114
rect 248690 151026 248870 151114
rect 248978 151026 249158 151114
rect 249266 151026 249446 151114
rect 249554 151026 249734 151114
rect 249842 151026 250022 151114
rect 250130 151026 250310 151114
rect 250564 151026 250744 151114
rect 360436 151026 360560 151114
rect 360814 151026 360994 151114
rect 361102 151026 361282 151114
rect 361390 151026 361570 151114
rect 361678 151026 361858 151114
rect 361966 151026 362146 151114
rect 362254 151026 362434 151114
rect 362542 151026 362722 151114
rect 362830 151026 363010 151114
rect 363264 151026 363444 151114
rect 363552 151026 363732 151114
rect 363840 151026 364020 151114
rect 364128 151026 364308 151114
rect 364416 151026 364596 151114
rect 364704 151026 364884 151114
rect 364992 151026 365172 151114
rect 365280 151026 365460 151114
rect 365714 151026 365894 151114
rect 366002 151026 366182 151114
rect 366290 151026 366470 151114
rect 366578 151026 366758 151114
rect 366866 151026 367046 151114
rect 367154 151026 367334 151114
rect 367442 151026 367622 151114
rect 367730 151026 367910 151114
rect 243214 150810 243394 150898
rect 243502 150810 243682 150898
rect 243790 150810 243970 150898
rect 244078 150810 244258 150898
rect 244366 150810 244546 150898
rect 244654 150810 244834 150898
rect 244942 150810 245122 150898
rect 245230 150810 245410 150898
rect 245664 150810 245844 150898
rect 245952 150810 246132 150898
rect 246240 150810 246420 150898
rect 246528 150810 246708 150898
rect 246816 150810 246996 150898
rect 247104 150810 247284 150898
rect 247392 150810 247572 150898
rect 247680 150810 247860 150898
rect 248114 150810 248294 150898
rect 248402 150810 248582 150898
rect 248690 150810 248870 150898
rect 248978 150810 249158 150898
rect 249266 150810 249446 150898
rect 249554 150810 249734 150898
rect 249842 150810 250022 150898
rect 250130 150810 250310 150898
rect 250564 150810 250744 150898
rect 360436 150810 360560 150898
rect 360814 150810 360994 150898
rect 361102 150810 361282 150898
rect 361390 150810 361570 150898
rect 361678 150810 361858 150898
rect 361966 150810 362146 150898
rect 362254 150810 362434 150898
rect 362542 150810 362722 150898
rect 362830 150810 363010 150898
rect 363264 150810 363444 150898
rect 363552 150810 363732 150898
rect 363840 150810 364020 150898
rect 364128 150810 364308 150898
rect 364416 150810 364596 150898
rect 364704 150810 364884 150898
rect 364992 150810 365172 150898
rect 365280 150810 365460 150898
rect 365714 150810 365894 150898
rect 366002 150810 366182 150898
rect 366290 150810 366470 150898
rect 366578 150810 366758 150898
rect 366866 150810 367046 150898
rect 367154 150810 367334 150898
rect 367442 150810 367622 150898
rect 367730 150810 367910 150898
rect 243214 150334 243394 150422
rect 243502 150334 243682 150422
rect 243790 150334 243970 150422
rect 244078 150334 244258 150422
rect 244366 150334 244546 150422
rect 244654 150334 244834 150422
rect 244942 150334 245122 150422
rect 245230 150334 245410 150422
rect 245664 150334 245844 150422
rect 245952 150334 246132 150422
rect 246240 150334 246420 150422
rect 246528 150334 246708 150422
rect 246816 150334 246996 150422
rect 247104 150334 247284 150422
rect 247392 150334 247572 150422
rect 247680 150334 247860 150422
rect 248114 150334 248294 150422
rect 248402 150334 248582 150422
rect 248690 150334 248870 150422
rect 248978 150334 249158 150422
rect 249266 150334 249446 150422
rect 249554 150334 249734 150422
rect 249842 150334 250022 150422
rect 250130 150334 250310 150422
rect 250564 150334 250744 150422
rect 360436 150364 360560 150422
rect 250852 150334 251032 150364
rect 251140 150334 251320 150364
rect 251428 150334 251608 150364
rect 251716 150334 251896 150364
rect 252004 150334 252184 150364
rect 252292 150334 252472 150364
rect 252580 150334 252760 150364
rect 253014 150334 253194 150364
rect 253302 150334 253482 150364
rect 253590 150334 253770 150364
rect 253878 150334 254058 150364
rect 254166 150334 254346 150364
rect 254454 150334 254634 150364
rect 254742 150334 254922 150364
rect 255030 150334 255210 150364
rect 255464 150334 255644 150364
rect 255752 150334 255932 150364
rect 256040 150334 256220 150364
rect 256328 150334 256508 150364
rect 256616 150334 256796 150364
rect 256904 150334 257084 150364
rect 257192 150334 257372 150364
rect 257480 150334 257660 150364
rect 257914 150334 258094 150364
rect 258202 150334 258382 150364
rect 258490 150334 258670 150364
rect 258778 150334 258958 150364
rect 259066 150334 259246 150364
rect 259354 150334 259534 150364
rect 259642 150334 259822 150364
rect 259930 150334 260110 150364
rect 260364 150334 260544 150364
rect 260652 150334 260832 150364
rect 260940 150334 261120 150364
rect 261228 150334 261408 150364
rect 261516 150334 261696 150364
rect 261804 150334 261984 150364
rect 262092 150334 262272 150364
rect 262380 150334 262560 150364
rect 262814 150334 262994 150364
rect 263102 150334 263282 150364
rect 263390 150334 263570 150364
rect 263678 150334 263858 150364
rect 263966 150334 264146 150364
rect 264254 150334 264434 150364
rect 264542 150334 264722 150364
rect 264830 150334 265010 150364
rect 265264 150334 265444 150364
rect 265552 150334 265732 150364
rect 265840 150334 266020 150364
rect 266128 150334 266308 150364
rect 266416 150334 266596 150364
rect 266704 150334 266884 150364
rect 266992 150334 267172 150364
rect 267280 150334 267460 150364
rect 267714 150334 267894 150364
rect 268002 150334 268182 150364
rect 268290 150334 268470 150364
rect 268578 150334 268758 150364
rect 268866 150334 269046 150364
rect 269154 150334 269334 150364
rect 269442 150334 269622 150364
rect 269730 150334 269910 150364
rect 270164 150334 270344 150364
rect 270452 150334 270632 150364
rect 270740 150334 270920 150364
rect 271028 150334 271208 150364
rect 271316 150334 271496 150364
rect 271604 150334 271784 150364
rect 271892 150334 272072 150364
rect 272180 150334 272360 150364
rect 272614 150334 272794 150364
rect 272902 150334 273082 150364
rect 273190 150334 273370 150364
rect 273478 150334 273658 150364
rect 273766 150334 273946 150364
rect 274054 150334 274234 150364
rect 274342 150334 274522 150364
rect 274630 150334 274810 150364
rect 275064 150334 275244 150364
rect 275352 150334 275532 150364
rect 275640 150334 275820 150364
rect 275928 150334 276108 150364
rect 276216 150334 276396 150364
rect 276504 150334 276684 150364
rect 276792 150334 276972 150364
rect 277080 150334 277260 150364
rect 277514 150334 277694 150364
rect 277802 150334 277982 150364
rect 278090 150334 278270 150364
rect 278378 150334 278558 150364
rect 278666 150334 278846 150364
rect 278954 150334 279134 150364
rect 279242 150334 279422 150364
rect 279530 150334 279710 150364
rect 279964 150334 280144 150364
rect 280252 150334 280432 150364
rect 280540 150334 280720 150364
rect 280828 150334 281008 150364
rect 281116 150334 281296 150364
rect 281404 150334 281584 150364
rect 281692 150334 281872 150364
rect 281980 150334 282160 150364
rect 282414 150334 282594 150364
rect 282702 150334 282882 150364
rect 282990 150334 283170 150364
rect 283278 150334 283458 150364
rect 283566 150334 283746 150364
rect 283854 150334 284034 150364
rect 284142 150334 284322 150364
rect 284430 150334 284610 150364
rect 284864 150334 285044 150364
rect 285152 150334 285332 150364
rect 285440 150334 285620 150364
rect 285728 150334 285908 150364
rect 286016 150334 286196 150364
rect 286304 150334 286484 150364
rect 286592 150334 286772 150364
rect 286880 150334 287060 150364
rect 287314 150334 287494 150364
rect 287602 150334 287782 150364
rect 287890 150334 288070 150364
rect 288178 150334 288358 150364
rect 288466 150334 288646 150364
rect 288754 150334 288934 150364
rect 289042 150334 289222 150364
rect 289330 150334 289510 150364
rect 289764 150334 289944 150364
rect 290052 150334 290232 150364
rect 290340 150334 290520 150364
rect 290628 150334 290808 150364
rect 290916 150334 291096 150364
rect 291204 150334 291384 150364
rect 291492 150334 291672 150364
rect 291780 150334 291960 150364
rect 292214 150334 292394 150364
rect 292502 150334 292682 150364
rect 292790 150334 292970 150364
rect 293078 150334 293258 150364
rect 293366 150334 293546 150364
rect 293654 150334 293834 150364
rect 293942 150334 294122 150364
rect 294230 150334 294410 150364
rect 294664 150334 294844 150364
rect 294952 150334 295132 150364
rect 295240 150334 295420 150364
rect 295528 150334 295708 150364
rect 295816 150334 295996 150364
rect 296104 150334 296284 150364
rect 296392 150334 296572 150364
rect 296680 150334 296860 150364
rect 297114 150334 297294 150364
rect 297402 150334 297582 150364
rect 297690 150334 297870 150364
rect 297978 150334 298158 150364
rect 298266 150334 298446 150364
rect 298554 150334 298734 150364
rect 298842 150334 299022 150364
rect 299130 150334 299310 150364
rect 299564 150334 299744 150364
rect 299852 150334 300032 150364
rect 300140 150334 300320 150364
rect 300428 150334 300608 150364
rect 300716 150334 300896 150364
rect 301004 150334 301184 150364
rect 301292 150334 301472 150364
rect 301580 150334 301760 150364
rect 302014 150334 302194 150364
rect 302302 150334 302482 150364
rect 302590 150334 302770 150364
rect 302878 150334 303058 150364
rect 303166 150334 303346 150364
rect 303454 150334 303634 150364
rect 303742 150334 303922 150364
rect 304030 150334 304210 150364
rect 304464 150334 304644 150364
rect 304752 150334 304932 150364
rect 305040 150334 305220 150364
rect 305328 150334 305508 150364
rect 305616 150334 305796 150364
rect 305904 150334 306084 150364
rect 306192 150334 306372 150364
rect 306480 150334 306660 150364
rect 306914 150334 307094 150364
rect 307202 150334 307382 150364
rect 307490 150334 307670 150364
rect 307778 150334 307958 150364
rect 308066 150334 308246 150364
rect 308354 150334 308534 150364
rect 308642 150334 308822 150364
rect 308930 150334 309110 150364
rect 309364 150334 309544 150364
rect 309652 150334 309832 150364
rect 309940 150334 310120 150364
rect 310228 150334 310408 150364
rect 310516 150334 310696 150364
rect 310804 150334 310984 150364
rect 311092 150334 311272 150364
rect 311380 150334 311560 150364
rect 311814 150334 311994 150364
rect 312102 150334 312282 150364
rect 312390 150334 312570 150364
rect 312678 150334 312858 150364
rect 312966 150334 313146 150364
rect 313254 150334 313434 150364
rect 313542 150334 313722 150364
rect 313830 150334 314010 150364
rect 314264 150334 314444 150364
rect 314552 150334 314732 150364
rect 314840 150334 315020 150364
rect 315128 150334 315308 150364
rect 315416 150334 315596 150364
rect 315704 150334 315884 150364
rect 315992 150334 316172 150364
rect 316280 150334 316460 150364
rect 316714 150334 316894 150364
rect 317002 150334 317182 150364
rect 317290 150334 317470 150364
rect 317578 150334 317758 150364
rect 317866 150334 318046 150364
rect 318154 150334 318334 150364
rect 318442 150334 318622 150364
rect 318730 150334 318910 150364
rect 319164 150334 319344 150364
rect 319452 150334 319632 150364
rect 319740 150334 319920 150364
rect 320028 150334 320208 150364
rect 320316 150334 320496 150364
rect 320604 150334 320784 150364
rect 320892 150334 321072 150364
rect 321180 150334 321360 150364
rect 321614 150334 321794 150364
rect 321902 150334 322082 150364
rect 322190 150334 322370 150364
rect 322478 150334 322658 150364
rect 322766 150334 322946 150364
rect 323054 150334 323234 150364
rect 323342 150334 323522 150364
rect 323630 150334 323810 150364
rect 324064 150334 324244 150364
rect 324352 150334 324532 150364
rect 324640 150334 324820 150364
rect 324928 150334 325108 150364
rect 325216 150334 325396 150364
rect 325504 150334 325684 150364
rect 325792 150334 325972 150364
rect 326080 150334 326260 150364
rect 326514 150334 326694 150364
rect 326802 150334 326982 150364
rect 327090 150334 327270 150364
rect 327378 150334 327558 150364
rect 327666 150334 327846 150364
rect 327954 150334 328134 150364
rect 328242 150334 328422 150364
rect 328530 150334 328710 150364
rect 328964 150334 329144 150364
rect 329252 150334 329432 150364
rect 329540 150334 329720 150364
rect 329828 150334 330008 150364
rect 330116 150334 330296 150364
rect 330404 150334 330584 150364
rect 330692 150334 330872 150364
rect 330980 150334 331160 150364
rect 331414 150334 331594 150364
rect 331702 150334 331882 150364
rect 331990 150334 332170 150364
rect 332278 150334 332458 150364
rect 332566 150334 332746 150364
rect 332854 150334 333034 150364
rect 333142 150334 333322 150364
rect 333430 150334 333610 150364
rect 333864 150334 334044 150364
rect 334152 150334 334332 150364
rect 334440 150334 334620 150364
rect 334728 150334 334908 150364
rect 335016 150334 335196 150364
rect 335304 150334 335484 150364
rect 335592 150334 335772 150364
rect 335880 150334 336060 150364
rect 336314 150334 336494 150364
rect 336602 150334 336782 150364
rect 336890 150334 337070 150364
rect 337178 150334 337358 150364
rect 337466 150334 337646 150364
rect 337754 150334 337934 150364
rect 338042 150334 338222 150364
rect 338330 150334 338510 150364
rect 338764 150334 338944 150364
rect 339052 150334 339232 150364
rect 339340 150334 339520 150364
rect 339628 150334 339808 150364
rect 339916 150334 340096 150364
rect 340204 150334 340384 150364
rect 340492 150334 340672 150364
rect 340780 150334 340960 150364
rect 341214 150334 341394 150364
rect 341502 150334 341682 150364
rect 341790 150334 341970 150364
rect 342078 150334 342258 150364
rect 342366 150334 342546 150364
rect 342654 150334 342834 150364
rect 342942 150334 343122 150364
rect 343230 150334 343410 150364
rect 343664 150334 343844 150364
rect 343952 150334 344132 150364
rect 344240 150334 344420 150364
rect 344528 150334 344708 150364
rect 344816 150334 344996 150364
rect 345104 150334 345284 150364
rect 345392 150334 345572 150364
rect 345680 150334 345860 150364
rect 346114 150334 346294 150364
rect 346402 150334 346582 150364
rect 346690 150334 346870 150364
rect 346978 150334 347158 150364
rect 347266 150334 347446 150364
rect 347554 150334 347734 150364
rect 347842 150334 348022 150364
rect 348130 150334 348310 150364
rect 348564 150334 348744 150364
rect 348852 150334 349032 150364
rect 349140 150334 349320 150364
rect 349428 150334 349608 150364
rect 349716 150334 349896 150364
rect 350004 150334 350184 150364
rect 350292 150334 350472 150364
rect 350580 150334 350760 150364
rect 351014 150334 351194 150364
rect 351302 150334 351482 150364
rect 351590 150334 351770 150364
rect 351878 150334 352058 150364
rect 352166 150334 352346 150364
rect 352454 150334 352634 150364
rect 352742 150334 352922 150364
rect 353030 150334 353210 150364
rect 353464 150334 353644 150364
rect 353752 150334 353932 150364
rect 354040 150334 354220 150364
rect 354328 150334 354508 150364
rect 354616 150334 354796 150364
rect 354904 150334 355084 150364
rect 355192 150334 355372 150364
rect 355480 150334 355660 150364
rect 355914 150334 356094 150364
rect 356202 150334 356382 150364
rect 356490 150334 356670 150364
rect 356778 150334 356958 150364
rect 357066 150334 357246 150364
rect 357354 150334 357534 150364
rect 357642 150334 357822 150364
rect 357930 150334 358110 150364
rect 358364 150334 358544 150364
rect 358652 150334 358832 150364
rect 358940 150334 359120 150364
rect 359228 150334 359408 150364
rect 359516 150334 359696 150364
rect 359804 150334 359984 150364
rect 360092 150334 360272 150364
rect 360380 150334 360560 150364
rect 360814 150334 360994 150422
rect 361102 150334 361282 150422
rect 361390 150334 361570 150422
rect 361678 150334 361858 150422
rect 361966 150334 362146 150422
rect 362254 150334 362434 150422
rect 362542 150334 362722 150422
rect 362830 150334 363010 150422
rect 363264 150334 363444 150422
rect 363552 150334 363732 150422
rect 363840 150334 364020 150422
rect 364128 150334 364308 150422
rect 364416 150334 364596 150422
rect 364704 150334 364884 150422
rect 364992 150334 365172 150422
rect 365280 150334 365460 150422
rect 365714 150334 365894 150422
rect 366002 150334 366182 150422
rect 366290 150334 366470 150422
rect 366578 150334 366758 150422
rect 366866 150334 367046 150422
rect 367154 150334 367334 150422
rect 367442 150334 367622 150422
rect 367730 150334 367910 150422
rect 243214 150118 243394 150206
rect 243502 150118 243682 150206
rect 243790 150118 243970 150206
rect 244078 150118 244258 150206
rect 244366 150118 244546 150206
rect 244654 150118 244834 150206
rect 244942 150118 245122 150206
rect 245230 150118 245410 150206
rect 245664 150118 245844 150206
rect 245952 150118 246132 150206
rect 246240 150118 246420 150206
rect 246528 150118 246708 150206
rect 246816 150118 246996 150206
rect 247104 150118 247284 150206
rect 247392 150118 247572 150206
rect 247680 150118 247860 150206
rect 248114 150118 248294 150206
rect 248402 150118 248582 150206
rect 248690 150118 248870 150206
rect 248978 150118 249158 150206
rect 249266 150118 249446 150206
rect 249554 150118 249734 150206
rect 249842 150118 250022 150206
rect 250130 150118 250310 150206
rect 250564 150118 250744 150206
rect 250852 150118 251032 150206
rect 251140 150118 251320 150206
rect 251428 150118 251608 150206
rect 251716 150118 251896 150206
rect 252004 150118 252184 150206
rect 252292 150118 252472 150206
rect 252580 150118 252760 150206
rect 253014 150118 253194 150206
rect 253302 150118 253482 150206
rect 253590 150118 253770 150206
rect 253878 150118 254058 150206
rect 254166 150118 254346 150206
rect 254454 150118 254634 150206
rect 254742 150118 254922 150206
rect 255030 150118 255210 150206
rect 255464 150118 255644 150206
rect 255752 150118 255932 150206
rect 256040 150118 256220 150206
rect 256328 150118 256508 150206
rect 256616 150118 256796 150206
rect 256904 150118 257084 150206
rect 257192 150118 257372 150206
rect 257480 150118 257660 150206
rect 257914 150118 258094 150206
rect 258202 150118 258382 150206
rect 258490 150118 258670 150206
rect 258778 150118 258958 150206
rect 259066 150118 259246 150206
rect 259354 150118 259534 150206
rect 259642 150118 259822 150206
rect 259930 150118 260110 150206
rect 260364 150118 260544 150206
rect 260652 150118 260832 150206
rect 260940 150118 261120 150206
rect 261228 150118 261408 150206
rect 261516 150118 261696 150206
rect 261804 150118 261984 150206
rect 262092 150118 262272 150206
rect 262380 150118 262560 150206
rect 262814 150118 262994 150206
rect 263102 150118 263282 150206
rect 263390 150118 263570 150206
rect 263678 150118 263858 150206
rect 263966 150118 264146 150206
rect 264254 150118 264434 150206
rect 264542 150118 264722 150206
rect 264830 150118 265010 150206
rect 265264 150118 265444 150206
rect 265552 150118 265732 150206
rect 265840 150118 266020 150206
rect 266128 150118 266308 150206
rect 266416 150118 266596 150206
rect 266704 150118 266884 150206
rect 266992 150118 267172 150206
rect 267280 150118 267460 150206
rect 267714 150118 267894 150206
rect 268002 150118 268182 150206
rect 268290 150118 268470 150206
rect 268578 150118 268758 150206
rect 268866 150118 269046 150206
rect 269154 150118 269334 150206
rect 269442 150118 269622 150206
rect 269730 150118 269910 150206
rect 270164 150118 270344 150206
rect 270452 150118 270632 150206
rect 270740 150118 270920 150206
rect 271028 150118 271208 150206
rect 271316 150118 271496 150206
rect 271604 150118 271784 150206
rect 271892 150118 272072 150206
rect 272180 150118 272360 150206
rect 272614 150118 272794 150206
rect 272902 150118 273082 150206
rect 273190 150118 273370 150206
rect 273478 150118 273658 150206
rect 273766 150118 273946 150206
rect 274054 150118 274234 150206
rect 274342 150118 274522 150206
rect 274630 150118 274810 150206
rect 275064 150118 275244 150206
rect 275352 150118 275532 150206
rect 275640 150118 275820 150206
rect 275928 150118 276108 150206
rect 276216 150118 276396 150206
rect 276504 150118 276684 150206
rect 276792 150118 276972 150206
rect 277080 150118 277260 150206
rect 277514 150118 277694 150206
rect 277802 150118 277982 150206
rect 278090 150118 278270 150206
rect 278378 150118 278558 150206
rect 278666 150118 278846 150206
rect 278954 150118 279134 150206
rect 279242 150118 279422 150206
rect 279530 150118 279710 150206
rect 279964 150118 280144 150206
rect 280252 150118 280432 150206
rect 280540 150118 280720 150206
rect 280828 150118 281008 150206
rect 281116 150118 281296 150206
rect 281404 150118 281584 150206
rect 281692 150118 281872 150206
rect 281980 150118 282160 150206
rect 282414 150118 282594 150206
rect 282702 150118 282882 150206
rect 282990 150118 283170 150206
rect 283278 150118 283458 150206
rect 283566 150118 283746 150206
rect 283854 150118 284034 150206
rect 284142 150118 284322 150206
rect 284430 150118 284610 150206
rect 284864 150118 285044 150206
rect 285152 150118 285332 150206
rect 285440 150118 285620 150206
rect 285728 150118 285908 150206
rect 286016 150118 286196 150206
rect 286304 150118 286484 150206
rect 286592 150118 286772 150206
rect 286880 150118 287060 150206
rect 287314 150118 287494 150206
rect 287602 150118 287782 150206
rect 287890 150118 288070 150206
rect 288178 150118 288358 150206
rect 288466 150118 288646 150206
rect 288754 150118 288934 150206
rect 289042 150118 289222 150206
rect 289330 150118 289510 150206
rect 289764 150118 289944 150206
rect 290052 150118 290232 150206
rect 290340 150118 290520 150206
rect 290628 150118 290808 150206
rect 290916 150118 291096 150206
rect 291204 150118 291384 150206
rect 291492 150118 291672 150206
rect 291780 150118 291960 150206
rect 292214 150118 292394 150206
rect 292502 150118 292682 150206
rect 292790 150118 292970 150206
rect 293078 150118 293258 150206
rect 293366 150118 293546 150206
rect 293654 150118 293834 150206
rect 293942 150118 294122 150206
rect 294230 150118 294410 150206
rect 294664 150118 294844 150206
rect 294952 150118 295132 150206
rect 295240 150118 295420 150206
rect 295528 150118 295708 150206
rect 295816 150118 295996 150206
rect 296104 150118 296284 150206
rect 296392 150118 296572 150206
rect 296680 150118 296860 150206
rect 297114 150118 297294 150206
rect 297402 150118 297582 150206
rect 297690 150118 297870 150206
rect 297978 150118 298158 150206
rect 298266 150118 298446 150206
rect 298554 150118 298734 150206
rect 298842 150118 299022 150206
rect 299130 150118 299310 150206
rect 299564 150118 299744 150206
rect 299852 150118 300032 150206
rect 300140 150118 300320 150206
rect 300428 150118 300608 150206
rect 300716 150118 300896 150206
rect 301004 150118 301184 150206
rect 301292 150118 301472 150206
rect 301580 150118 301760 150206
rect 302014 150118 302194 150206
rect 302302 150118 302482 150206
rect 302590 150118 302770 150206
rect 302878 150118 303058 150206
rect 303166 150118 303346 150206
rect 303454 150118 303634 150206
rect 303742 150118 303922 150206
rect 304030 150118 304210 150206
rect 304464 150118 304644 150206
rect 304752 150118 304932 150206
rect 305040 150118 305220 150206
rect 305328 150118 305508 150206
rect 305616 150118 305796 150206
rect 305904 150118 306084 150206
rect 306192 150118 306372 150206
rect 306480 150118 306660 150206
rect 306914 150118 307094 150206
rect 307202 150118 307382 150206
rect 307490 150118 307670 150206
rect 307778 150118 307958 150206
rect 308066 150118 308246 150206
rect 308354 150118 308534 150206
rect 308642 150118 308822 150206
rect 308930 150118 309110 150206
rect 309364 150118 309544 150206
rect 309652 150118 309832 150206
rect 309940 150118 310120 150206
rect 310228 150118 310408 150206
rect 310516 150118 310696 150206
rect 310804 150118 310984 150206
rect 311092 150118 311272 150206
rect 311380 150118 311560 150206
rect 311814 150118 311994 150206
rect 312102 150118 312282 150206
rect 312390 150118 312570 150206
rect 312678 150118 312858 150206
rect 312966 150118 313146 150206
rect 313254 150118 313434 150206
rect 313542 150118 313722 150206
rect 313830 150118 314010 150206
rect 314264 150118 314444 150206
rect 314552 150118 314732 150206
rect 314840 150118 315020 150206
rect 315128 150118 315308 150206
rect 315416 150118 315596 150206
rect 315704 150118 315884 150206
rect 315992 150118 316172 150206
rect 316280 150118 316460 150206
rect 316714 150118 316894 150206
rect 317002 150118 317182 150206
rect 317290 150118 317470 150206
rect 317578 150118 317758 150206
rect 317866 150118 318046 150206
rect 318154 150118 318334 150206
rect 318442 150118 318622 150206
rect 318730 150118 318910 150206
rect 319164 150118 319344 150206
rect 319452 150118 319632 150206
rect 319740 150118 319920 150206
rect 320028 150118 320208 150206
rect 320316 150118 320496 150206
rect 320604 150118 320784 150206
rect 320892 150118 321072 150206
rect 321180 150118 321360 150206
rect 321614 150118 321794 150206
rect 321902 150118 322082 150206
rect 322190 150118 322370 150206
rect 322478 150118 322658 150206
rect 322766 150118 322946 150206
rect 323054 150118 323234 150206
rect 323342 150118 323522 150206
rect 323630 150118 323810 150206
rect 324064 150118 324244 150206
rect 324352 150118 324532 150206
rect 324640 150118 324820 150206
rect 324928 150118 325108 150206
rect 325216 150118 325396 150206
rect 325504 150118 325684 150206
rect 325792 150118 325972 150206
rect 326080 150118 326260 150206
rect 326514 150118 326694 150206
rect 326802 150118 326982 150206
rect 327090 150118 327270 150206
rect 327378 150118 327558 150206
rect 327666 150118 327846 150206
rect 327954 150118 328134 150206
rect 328242 150118 328422 150206
rect 328530 150118 328710 150206
rect 328964 150118 329144 150206
rect 329252 150118 329432 150206
rect 329540 150118 329720 150206
rect 329828 150118 330008 150206
rect 330116 150118 330296 150206
rect 330404 150118 330584 150206
rect 330692 150118 330872 150206
rect 330980 150118 331160 150206
rect 331414 150118 331594 150206
rect 331702 150118 331882 150206
rect 331990 150118 332170 150206
rect 332278 150118 332458 150206
rect 332566 150118 332746 150206
rect 332854 150118 333034 150206
rect 333142 150118 333322 150206
rect 333430 150118 333610 150206
rect 333864 150118 334044 150206
rect 334152 150118 334332 150206
rect 334440 150118 334620 150206
rect 334728 150118 334908 150206
rect 335016 150118 335196 150206
rect 335304 150118 335484 150206
rect 335592 150118 335772 150206
rect 335880 150118 336060 150206
rect 336314 150118 336494 150206
rect 336602 150118 336782 150206
rect 336890 150118 337070 150206
rect 337178 150118 337358 150206
rect 337466 150118 337646 150206
rect 337754 150118 337934 150206
rect 338042 150118 338222 150206
rect 338330 150118 338510 150206
rect 338764 150118 338944 150206
rect 339052 150118 339232 150206
rect 339340 150118 339520 150206
rect 339628 150118 339808 150206
rect 339916 150118 340096 150206
rect 340204 150118 340384 150206
rect 340492 150118 340672 150206
rect 340780 150118 340960 150206
rect 341214 150118 341394 150206
rect 341502 150118 341682 150206
rect 341790 150118 341970 150206
rect 342078 150118 342258 150206
rect 342366 150118 342546 150206
rect 342654 150118 342834 150206
rect 342942 150118 343122 150206
rect 343230 150118 343410 150206
rect 343664 150118 343844 150206
rect 343952 150118 344132 150206
rect 344240 150118 344420 150206
rect 344528 150118 344708 150206
rect 344816 150118 344996 150206
rect 345104 150118 345284 150206
rect 345392 150118 345572 150206
rect 345680 150118 345860 150206
rect 346114 150118 346294 150206
rect 346402 150118 346582 150206
rect 346690 150118 346870 150206
rect 346978 150118 347158 150206
rect 347266 150118 347446 150206
rect 347554 150118 347734 150206
rect 347842 150118 348022 150206
rect 348130 150118 348310 150206
rect 348564 150118 348744 150206
rect 348852 150118 349032 150206
rect 349140 150118 349320 150206
rect 349428 150118 349608 150206
rect 349716 150118 349896 150206
rect 350004 150118 350184 150206
rect 350292 150118 350472 150206
rect 350580 150118 350760 150206
rect 351014 150118 351194 150206
rect 351302 150118 351482 150206
rect 351590 150118 351770 150206
rect 351878 150118 352058 150206
rect 352166 150118 352346 150206
rect 352454 150118 352634 150206
rect 352742 150118 352922 150206
rect 353030 150118 353210 150206
rect 353464 150118 353644 150206
rect 353752 150118 353932 150206
rect 354040 150118 354220 150206
rect 354328 150118 354508 150206
rect 354616 150118 354796 150206
rect 354904 150118 355084 150206
rect 355192 150118 355372 150206
rect 355480 150118 355660 150206
rect 355914 150118 356094 150206
rect 356202 150118 356382 150206
rect 356490 150118 356670 150206
rect 356778 150118 356958 150206
rect 357066 150118 357246 150206
rect 357354 150118 357534 150206
rect 357642 150118 357822 150206
rect 357930 150118 358110 150206
rect 358364 150118 358544 150206
rect 358652 150118 358832 150206
rect 358940 150118 359120 150206
rect 359228 150118 359408 150206
rect 359516 150118 359696 150206
rect 359804 150118 359984 150206
rect 360092 150118 360272 150206
rect 360380 150118 360560 150206
rect 360814 150118 360994 150206
rect 361102 150118 361282 150206
rect 361390 150118 361570 150206
rect 361678 150118 361858 150206
rect 361966 150118 362146 150206
rect 362254 150118 362434 150206
rect 362542 150118 362722 150206
rect 362830 150118 363010 150206
rect 363264 150118 363444 150206
rect 363552 150118 363732 150206
rect 363840 150118 364020 150206
rect 364128 150118 364308 150206
rect 364416 150118 364596 150206
rect 364704 150118 364884 150206
rect 364992 150118 365172 150206
rect 365280 150118 365460 150206
rect 365714 150118 365894 150206
rect 366002 150118 366182 150206
rect 366290 150118 366470 150206
rect 366578 150118 366758 150206
rect 366866 150118 367046 150206
rect 367154 150118 367334 150206
rect 367442 150118 367622 150206
rect 367730 150118 367910 150206
rect 243214 149642 243394 149730
rect 243502 149642 243682 149730
rect 243790 149642 243970 149730
rect 244078 149642 244258 149730
rect 244366 149642 244546 149730
rect 244654 149642 244834 149730
rect 244942 149642 245122 149730
rect 245230 149642 245410 149730
rect 245664 149642 245844 149730
rect 245952 149642 246132 149730
rect 246240 149642 246420 149730
rect 246528 149642 246708 149730
rect 246816 149642 246996 149730
rect 247104 149642 247284 149730
rect 247392 149642 247572 149730
rect 247680 149642 247860 149730
rect 248114 149642 248294 149730
rect 248402 149642 248582 149730
rect 248690 149642 248870 149730
rect 248978 149642 249158 149730
rect 249266 149642 249446 149730
rect 249554 149642 249734 149730
rect 249842 149642 250022 149730
rect 250130 149642 250310 149730
rect 250564 149642 250744 149730
rect 250852 149642 251032 149730
rect 251140 149642 251320 149730
rect 251428 149642 251608 149730
rect 251716 149642 251896 149730
rect 252004 149642 252184 149730
rect 252292 149642 252472 149730
rect 252580 149642 252760 149730
rect 253014 149642 253194 149730
rect 253302 149642 253482 149730
rect 253590 149642 253770 149730
rect 253878 149642 254058 149730
rect 254166 149642 254346 149730
rect 254454 149642 254634 149730
rect 254742 149642 254922 149730
rect 255030 149642 255210 149730
rect 255464 149642 255644 149730
rect 255752 149642 255932 149730
rect 256040 149642 256220 149730
rect 256328 149642 256508 149730
rect 256616 149642 256796 149730
rect 256904 149642 257084 149730
rect 257192 149642 257372 149730
rect 257480 149642 257660 149730
rect 257914 149642 258094 149730
rect 258202 149642 258382 149730
rect 258490 149642 258670 149730
rect 258778 149642 258958 149730
rect 259066 149642 259246 149730
rect 259354 149642 259534 149730
rect 259642 149642 259822 149730
rect 259930 149642 260110 149730
rect 260364 149642 260544 149730
rect 260652 149642 260832 149730
rect 260940 149642 261120 149730
rect 261228 149642 261408 149730
rect 261516 149642 261696 149730
rect 261804 149642 261984 149730
rect 262092 149642 262272 149730
rect 262380 149642 262560 149730
rect 262814 149642 262994 149730
rect 263102 149642 263282 149730
rect 263390 149642 263570 149730
rect 263678 149642 263858 149730
rect 263966 149642 264146 149730
rect 264254 149642 264434 149730
rect 264542 149642 264722 149730
rect 264830 149642 265010 149730
rect 265264 149642 265444 149730
rect 265552 149642 265732 149730
rect 265840 149642 266020 149730
rect 266128 149642 266308 149730
rect 266416 149642 266596 149730
rect 266704 149642 266884 149730
rect 266992 149642 267172 149730
rect 267280 149642 267460 149730
rect 267714 149642 267894 149730
rect 268002 149642 268182 149730
rect 268290 149642 268470 149730
rect 268578 149642 268758 149730
rect 268866 149642 269046 149730
rect 269154 149642 269334 149730
rect 269442 149642 269622 149730
rect 269730 149642 269910 149730
rect 270164 149642 270344 149730
rect 270452 149642 270632 149730
rect 270740 149642 270920 149730
rect 271028 149642 271208 149730
rect 271316 149642 271496 149730
rect 271604 149642 271784 149730
rect 271892 149642 272072 149730
rect 272180 149642 272360 149730
rect 272614 149642 272794 149730
rect 272902 149642 273082 149730
rect 273190 149642 273370 149730
rect 273478 149642 273658 149730
rect 273766 149642 273946 149730
rect 274054 149642 274234 149730
rect 274342 149642 274522 149730
rect 274630 149642 274810 149730
rect 275064 149642 275244 149730
rect 275352 149642 275532 149730
rect 275640 149642 275820 149730
rect 275928 149642 276108 149730
rect 276216 149642 276396 149730
rect 276504 149642 276684 149730
rect 276792 149642 276972 149730
rect 277080 149642 277260 149730
rect 277514 149642 277694 149730
rect 277802 149642 277982 149730
rect 278090 149642 278270 149730
rect 278378 149642 278558 149730
rect 278666 149642 278846 149730
rect 278954 149642 279134 149730
rect 279242 149642 279422 149730
rect 279530 149642 279710 149730
rect 279964 149642 280144 149730
rect 280252 149642 280432 149730
rect 280540 149642 280720 149730
rect 280828 149642 281008 149730
rect 281116 149642 281296 149730
rect 281404 149642 281584 149730
rect 281692 149642 281872 149730
rect 281980 149642 282160 149730
rect 282414 149642 282594 149730
rect 282702 149642 282882 149730
rect 282990 149642 283170 149730
rect 283278 149642 283458 149730
rect 283566 149642 283746 149730
rect 283854 149642 284034 149730
rect 284142 149642 284322 149730
rect 284430 149642 284610 149730
rect 284864 149642 285044 149730
rect 285152 149642 285332 149730
rect 285440 149642 285620 149730
rect 285728 149642 285908 149730
rect 286016 149642 286196 149730
rect 286304 149642 286484 149730
rect 286592 149642 286772 149730
rect 286880 149642 287060 149730
rect 287314 149642 287494 149730
rect 287602 149642 287782 149730
rect 287890 149642 288070 149730
rect 288178 149642 288358 149730
rect 288466 149642 288646 149730
rect 288754 149642 288934 149730
rect 289042 149642 289222 149730
rect 289330 149642 289510 149730
rect 289764 149642 289944 149730
rect 290052 149642 290232 149730
rect 290340 149642 290520 149730
rect 290628 149642 290808 149730
rect 290916 149642 291096 149730
rect 291204 149642 291384 149730
rect 291492 149642 291672 149730
rect 291780 149642 291960 149730
rect 292214 149642 292394 149730
rect 292502 149642 292682 149730
rect 292790 149642 292970 149730
rect 293078 149642 293258 149730
rect 293366 149642 293546 149730
rect 293654 149642 293834 149730
rect 293942 149642 294122 149730
rect 294230 149642 294410 149730
rect 294664 149642 294844 149730
rect 294952 149642 295132 149730
rect 295240 149642 295420 149730
rect 295528 149642 295708 149730
rect 295816 149642 295996 149730
rect 296104 149642 296284 149730
rect 296392 149642 296572 149730
rect 296680 149642 296860 149730
rect 297114 149642 297294 149730
rect 297402 149642 297582 149730
rect 297690 149642 297870 149730
rect 297978 149642 298158 149730
rect 298266 149642 298446 149730
rect 298554 149642 298734 149730
rect 298842 149642 299022 149730
rect 299130 149642 299310 149730
rect 299564 149642 299744 149730
rect 299852 149642 300032 149730
rect 300140 149642 300320 149730
rect 300428 149642 300608 149730
rect 300716 149642 300896 149730
rect 301004 149642 301184 149730
rect 301292 149642 301472 149730
rect 301580 149642 301760 149730
rect 302014 149642 302194 149730
rect 302302 149642 302482 149730
rect 302590 149642 302770 149730
rect 302878 149642 303058 149730
rect 303166 149642 303346 149730
rect 303454 149642 303634 149730
rect 303742 149642 303922 149730
rect 304030 149642 304210 149730
rect 304464 149642 304644 149730
rect 304752 149642 304932 149730
rect 305040 149642 305220 149730
rect 305328 149642 305508 149730
rect 305616 149642 305796 149730
rect 305904 149642 306084 149730
rect 306192 149642 306372 149730
rect 306480 149642 306660 149730
rect 306914 149642 307094 149730
rect 307202 149642 307382 149730
rect 307490 149642 307670 149730
rect 307778 149642 307958 149730
rect 308066 149642 308246 149730
rect 308354 149642 308534 149730
rect 308642 149642 308822 149730
rect 308930 149642 309110 149730
rect 309364 149642 309544 149730
rect 309652 149642 309832 149730
rect 309940 149642 310120 149730
rect 310228 149642 310408 149730
rect 310516 149642 310696 149730
rect 310804 149642 310984 149730
rect 311092 149642 311272 149730
rect 311380 149642 311560 149730
rect 311814 149642 311994 149730
rect 312102 149642 312282 149730
rect 312390 149642 312570 149730
rect 312678 149642 312858 149730
rect 312966 149642 313146 149730
rect 313254 149642 313434 149730
rect 313542 149642 313722 149730
rect 313830 149642 314010 149730
rect 314264 149642 314444 149730
rect 314552 149642 314732 149730
rect 314840 149642 315020 149730
rect 315128 149642 315308 149730
rect 315416 149642 315596 149730
rect 315704 149642 315884 149730
rect 315992 149642 316172 149730
rect 316280 149642 316460 149730
rect 316714 149642 316894 149730
rect 317002 149642 317182 149730
rect 317290 149642 317470 149730
rect 317578 149642 317758 149730
rect 317866 149642 318046 149730
rect 318154 149642 318334 149730
rect 318442 149642 318622 149730
rect 318730 149642 318910 149730
rect 319164 149642 319344 149730
rect 319452 149642 319632 149730
rect 319740 149642 319920 149730
rect 320028 149642 320208 149730
rect 320316 149642 320496 149730
rect 320604 149642 320784 149730
rect 320892 149642 321072 149730
rect 321180 149642 321360 149730
rect 321614 149642 321794 149730
rect 321902 149642 322082 149730
rect 322190 149642 322370 149730
rect 322478 149642 322658 149730
rect 322766 149642 322946 149730
rect 323054 149642 323234 149730
rect 323342 149642 323522 149730
rect 323630 149642 323810 149730
rect 324064 149642 324244 149730
rect 324352 149642 324532 149730
rect 324640 149642 324820 149730
rect 324928 149642 325108 149730
rect 325216 149642 325396 149730
rect 325504 149642 325684 149730
rect 325792 149642 325972 149730
rect 326080 149642 326260 149730
rect 326514 149642 326694 149730
rect 326802 149642 326982 149730
rect 327090 149642 327270 149730
rect 327378 149642 327558 149730
rect 327666 149642 327846 149730
rect 327954 149642 328134 149730
rect 328242 149642 328422 149730
rect 328530 149642 328710 149730
rect 328964 149642 329144 149730
rect 329252 149642 329432 149730
rect 329540 149642 329720 149730
rect 329828 149642 330008 149730
rect 330116 149642 330296 149730
rect 330404 149642 330584 149730
rect 330692 149642 330872 149730
rect 330980 149642 331160 149730
rect 331414 149642 331594 149730
rect 331702 149642 331882 149730
rect 331990 149642 332170 149730
rect 332278 149642 332458 149730
rect 332566 149642 332746 149730
rect 332854 149642 333034 149730
rect 333142 149642 333322 149730
rect 333430 149642 333610 149730
rect 333864 149642 334044 149730
rect 334152 149642 334332 149730
rect 334440 149642 334620 149730
rect 334728 149642 334908 149730
rect 335016 149642 335196 149730
rect 335304 149642 335484 149730
rect 335592 149642 335772 149730
rect 335880 149642 336060 149730
rect 336314 149642 336494 149730
rect 336602 149642 336782 149730
rect 336890 149642 337070 149730
rect 337178 149642 337358 149730
rect 337466 149642 337646 149730
rect 337754 149642 337934 149730
rect 338042 149642 338222 149730
rect 338330 149642 338510 149730
rect 338764 149642 338944 149730
rect 339052 149642 339232 149730
rect 339340 149642 339520 149730
rect 339628 149642 339808 149730
rect 339916 149642 340096 149730
rect 340204 149642 340384 149730
rect 340492 149642 340672 149730
rect 340780 149642 340960 149730
rect 341214 149642 341394 149730
rect 341502 149642 341682 149730
rect 341790 149642 341970 149730
rect 342078 149642 342258 149730
rect 342366 149642 342546 149730
rect 342654 149642 342834 149730
rect 342942 149642 343122 149730
rect 343230 149642 343410 149730
rect 343664 149642 343844 149730
rect 343952 149642 344132 149730
rect 344240 149642 344420 149730
rect 344528 149642 344708 149730
rect 344816 149642 344996 149730
rect 345104 149642 345284 149730
rect 345392 149642 345572 149730
rect 345680 149642 345860 149730
rect 346114 149642 346294 149730
rect 346402 149642 346582 149730
rect 346690 149642 346870 149730
rect 346978 149642 347158 149730
rect 347266 149642 347446 149730
rect 347554 149642 347734 149730
rect 347842 149642 348022 149730
rect 348130 149642 348310 149730
rect 348564 149642 348744 149730
rect 348852 149642 349032 149730
rect 349140 149642 349320 149730
rect 349428 149642 349608 149730
rect 349716 149642 349896 149730
rect 350004 149642 350184 149730
rect 350292 149642 350472 149730
rect 350580 149642 350760 149730
rect 351014 149642 351194 149730
rect 351302 149642 351482 149730
rect 351590 149642 351770 149730
rect 351878 149642 352058 149730
rect 352166 149642 352346 149730
rect 352454 149642 352634 149730
rect 352742 149642 352922 149730
rect 353030 149642 353210 149730
rect 353464 149642 353644 149730
rect 353752 149642 353932 149730
rect 354040 149642 354220 149730
rect 354328 149642 354508 149730
rect 354616 149642 354796 149730
rect 354904 149642 355084 149730
rect 355192 149642 355372 149730
rect 355480 149642 355660 149730
rect 355914 149642 356094 149730
rect 356202 149642 356382 149730
rect 356490 149642 356670 149730
rect 356778 149642 356958 149730
rect 357066 149642 357246 149730
rect 357354 149642 357534 149730
rect 357642 149642 357822 149730
rect 357930 149642 358110 149730
rect 358364 149642 358544 149730
rect 358652 149642 358832 149730
rect 358940 149642 359120 149730
rect 359228 149642 359408 149730
rect 359516 149642 359696 149730
rect 359804 149642 359984 149730
rect 360092 149642 360272 149730
rect 360380 149642 360560 149730
rect 360814 149642 360994 149730
rect 361102 149642 361282 149730
rect 361390 149642 361570 149730
rect 361678 149642 361858 149730
rect 361966 149642 362146 149730
rect 362254 149642 362434 149730
rect 362542 149642 362722 149730
rect 362830 149642 363010 149730
rect 363264 149642 363444 149730
rect 363552 149642 363732 149730
rect 363840 149642 364020 149730
rect 364128 149642 364308 149730
rect 364416 149642 364596 149730
rect 364704 149642 364884 149730
rect 364992 149642 365172 149730
rect 365280 149642 365460 149730
rect 365714 149642 365894 149730
rect 366002 149642 366182 149730
rect 366290 149642 366470 149730
rect 366578 149642 366758 149730
rect 366866 149642 367046 149730
rect 367154 149642 367334 149730
rect 367442 149642 367622 149730
rect 367730 149642 367910 149730
rect 243214 149426 243394 149514
rect 243502 149426 243682 149514
rect 243790 149426 243970 149514
rect 244078 149426 244258 149514
rect 244366 149426 244546 149514
rect 244654 149426 244834 149514
rect 244942 149426 245122 149514
rect 245230 149426 245410 149514
rect 245664 149426 245844 149514
rect 245952 149426 246132 149514
rect 246240 149426 246420 149514
rect 246528 149426 246708 149514
rect 246816 149426 246996 149514
rect 247104 149426 247284 149514
rect 247392 149426 247572 149514
rect 247680 149426 247860 149514
rect 248114 149426 248294 149514
rect 248402 149426 248582 149514
rect 248690 149426 248870 149514
rect 248978 149426 249158 149514
rect 249266 149426 249446 149514
rect 249554 149426 249734 149514
rect 249842 149426 250022 149514
rect 250130 149426 250310 149514
rect 250564 149426 250744 149514
rect 250852 149426 251032 149514
rect 251140 149426 251320 149514
rect 251428 149426 251608 149514
rect 251716 149426 251896 149514
rect 252004 149426 252184 149514
rect 252292 149426 252472 149514
rect 252580 149426 252760 149514
rect 253014 149426 253194 149514
rect 253302 149426 253482 149514
rect 253590 149426 253770 149514
rect 253878 149426 254058 149514
rect 254166 149426 254346 149514
rect 254454 149426 254634 149514
rect 254742 149426 254922 149514
rect 255030 149426 255210 149514
rect 255464 149426 255644 149514
rect 255752 149426 255932 149514
rect 256040 149426 256220 149514
rect 256328 149426 256508 149514
rect 256616 149426 256796 149514
rect 256904 149426 257084 149514
rect 257192 149426 257372 149514
rect 257480 149426 257660 149514
rect 257914 149426 258094 149514
rect 258202 149426 258382 149514
rect 258490 149426 258670 149514
rect 258778 149426 258958 149514
rect 259066 149426 259246 149514
rect 259354 149426 259534 149514
rect 259642 149426 259822 149514
rect 259930 149426 260110 149514
rect 260364 149426 260544 149514
rect 260652 149426 260832 149514
rect 260940 149426 261120 149514
rect 261228 149426 261408 149514
rect 261516 149426 261696 149514
rect 261804 149426 261984 149514
rect 262092 149426 262272 149514
rect 262380 149426 262560 149514
rect 262814 149426 262994 149514
rect 263102 149426 263282 149514
rect 263390 149426 263570 149514
rect 263678 149426 263858 149514
rect 263966 149426 264146 149514
rect 264254 149426 264434 149514
rect 264542 149426 264722 149514
rect 264830 149426 265010 149514
rect 265264 149426 265444 149514
rect 265552 149426 265732 149514
rect 265840 149426 266020 149514
rect 266128 149426 266308 149514
rect 266416 149426 266596 149514
rect 266704 149426 266884 149514
rect 266992 149426 267172 149514
rect 267280 149426 267460 149514
rect 267714 149426 267894 149514
rect 268002 149426 268182 149514
rect 268290 149426 268470 149514
rect 268578 149426 268758 149514
rect 268866 149426 269046 149514
rect 269154 149426 269334 149514
rect 269442 149426 269622 149514
rect 269730 149426 269910 149514
rect 270164 149426 270344 149514
rect 270452 149426 270632 149514
rect 270740 149426 270920 149514
rect 271028 149426 271208 149514
rect 271316 149426 271496 149514
rect 271604 149426 271784 149514
rect 271892 149426 272072 149514
rect 272180 149426 272360 149514
rect 272614 149426 272794 149514
rect 272902 149426 273082 149514
rect 273190 149426 273370 149514
rect 273478 149426 273658 149514
rect 273766 149426 273946 149514
rect 274054 149426 274234 149514
rect 274342 149426 274522 149514
rect 274630 149426 274810 149514
rect 275064 149426 275244 149514
rect 275352 149426 275532 149514
rect 275640 149426 275820 149514
rect 275928 149426 276108 149514
rect 276216 149426 276396 149514
rect 276504 149426 276684 149514
rect 276792 149426 276972 149514
rect 277080 149426 277260 149514
rect 277514 149426 277694 149514
rect 277802 149426 277982 149514
rect 278090 149426 278270 149514
rect 278378 149426 278558 149514
rect 278666 149426 278846 149514
rect 278954 149426 279134 149514
rect 279242 149426 279422 149514
rect 279530 149426 279710 149514
rect 279964 149426 280144 149514
rect 280252 149426 280432 149514
rect 280540 149426 280720 149514
rect 280828 149426 281008 149514
rect 281116 149426 281296 149514
rect 281404 149426 281584 149514
rect 281692 149426 281872 149514
rect 281980 149426 282160 149514
rect 282414 149426 282594 149514
rect 282702 149426 282882 149514
rect 282990 149426 283170 149514
rect 283278 149426 283458 149514
rect 283566 149426 283746 149514
rect 283854 149426 284034 149514
rect 284142 149426 284322 149514
rect 284430 149426 284610 149514
rect 284864 149426 285044 149514
rect 285152 149426 285332 149514
rect 285440 149426 285620 149514
rect 285728 149426 285908 149514
rect 286016 149426 286196 149514
rect 286304 149426 286484 149514
rect 286592 149426 286772 149514
rect 286880 149426 287060 149514
rect 287314 149426 287494 149514
rect 287602 149426 287782 149514
rect 287890 149426 288070 149514
rect 288178 149426 288358 149514
rect 288466 149426 288646 149514
rect 288754 149426 288934 149514
rect 289042 149426 289222 149514
rect 289330 149426 289510 149514
rect 289764 149426 289944 149514
rect 290052 149426 290232 149514
rect 290340 149426 290520 149514
rect 290628 149426 290808 149514
rect 290916 149426 291096 149514
rect 291204 149426 291384 149514
rect 291492 149426 291672 149514
rect 291780 149426 291960 149514
rect 292214 149426 292394 149514
rect 292502 149426 292682 149514
rect 292790 149426 292970 149514
rect 293078 149426 293258 149514
rect 293366 149426 293546 149514
rect 293654 149426 293834 149514
rect 293942 149426 294122 149514
rect 294230 149426 294410 149514
rect 294664 149426 294844 149514
rect 294952 149426 295132 149514
rect 295240 149426 295420 149514
rect 295528 149426 295708 149514
rect 295816 149426 295996 149514
rect 296104 149426 296284 149514
rect 296392 149426 296572 149514
rect 296680 149426 296860 149514
rect 297114 149426 297294 149514
rect 297402 149426 297582 149514
rect 297690 149426 297870 149514
rect 297978 149426 298158 149514
rect 298266 149426 298446 149514
rect 298554 149426 298734 149514
rect 298842 149426 299022 149514
rect 299130 149426 299310 149514
rect 299564 149426 299744 149514
rect 299852 149426 300032 149514
rect 300140 149426 300320 149514
rect 300428 149426 300608 149514
rect 300716 149426 300896 149514
rect 301004 149426 301184 149514
rect 301292 149426 301472 149514
rect 301580 149426 301760 149514
rect 302014 149426 302194 149514
rect 302302 149426 302482 149514
rect 302590 149426 302770 149514
rect 302878 149426 303058 149514
rect 303166 149426 303346 149514
rect 303454 149426 303634 149514
rect 303742 149426 303922 149514
rect 304030 149426 304210 149514
rect 304464 149426 304644 149514
rect 304752 149426 304932 149514
rect 305040 149426 305220 149514
rect 305328 149426 305508 149514
rect 305616 149426 305796 149514
rect 305904 149426 306084 149514
rect 306192 149426 306372 149514
rect 306480 149426 306660 149514
rect 306914 149426 307094 149514
rect 307202 149426 307382 149514
rect 307490 149426 307670 149514
rect 307778 149426 307958 149514
rect 308066 149426 308246 149514
rect 308354 149426 308534 149514
rect 308642 149426 308822 149514
rect 308930 149426 309110 149514
rect 309364 149426 309544 149514
rect 309652 149426 309832 149514
rect 309940 149426 310120 149514
rect 310228 149426 310408 149514
rect 310516 149426 310696 149514
rect 310804 149426 310984 149514
rect 311092 149426 311272 149514
rect 311380 149426 311560 149514
rect 311814 149426 311994 149514
rect 312102 149426 312282 149514
rect 312390 149426 312570 149514
rect 312678 149426 312858 149514
rect 312966 149426 313146 149514
rect 313254 149426 313434 149514
rect 313542 149426 313722 149514
rect 313830 149426 314010 149514
rect 314264 149426 314444 149514
rect 314552 149426 314732 149514
rect 314840 149426 315020 149514
rect 315128 149426 315308 149514
rect 315416 149426 315596 149514
rect 315704 149426 315884 149514
rect 315992 149426 316172 149514
rect 316280 149426 316460 149514
rect 316714 149426 316894 149514
rect 317002 149426 317182 149514
rect 317290 149426 317470 149514
rect 317578 149426 317758 149514
rect 317866 149426 318046 149514
rect 318154 149426 318334 149514
rect 318442 149426 318622 149514
rect 318730 149426 318910 149514
rect 319164 149426 319344 149514
rect 319452 149426 319632 149514
rect 319740 149426 319920 149514
rect 320028 149426 320208 149514
rect 320316 149426 320496 149514
rect 320604 149426 320784 149514
rect 320892 149426 321072 149514
rect 321180 149426 321360 149514
rect 321614 149426 321794 149514
rect 321902 149426 322082 149514
rect 322190 149426 322370 149514
rect 322478 149426 322658 149514
rect 322766 149426 322946 149514
rect 323054 149426 323234 149514
rect 323342 149426 323522 149514
rect 323630 149426 323810 149514
rect 324064 149426 324244 149514
rect 324352 149426 324532 149514
rect 324640 149426 324820 149514
rect 324928 149426 325108 149514
rect 325216 149426 325396 149514
rect 325504 149426 325684 149514
rect 325792 149426 325972 149514
rect 326080 149426 326260 149514
rect 326514 149426 326694 149514
rect 326802 149426 326982 149514
rect 327090 149426 327270 149514
rect 327378 149426 327558 149514
rect 327666 149426 327846 149514
rect 327954 149426 328134 149514
rect 328242 149426 328422 149514
rect 328530 149426 328710 149514
rect 328964 149426 329144 149514
rect 329252 149426 329432 149514
rect 329540 149426 329720 149514
rect 329828 149426 330008 149514
rect 330116 149426 330296 149514
rect 330404 149426 330584 149514
rect 330692 149426 330872 149514
rect 330980 149426 331160 149514
rect 331414 149426 331594 149514
rect 331702 149426 331882 149514
rect 331990 149426 332170 149514
rect 332278 149426 332458 149514
rect 332566 149426 332746 149514
rect 332854 149426 333034 149514
rect 333142 149426 333322 149514
rect 333430 149426 333610 149514
rect 333864 149426 334044 149514
rect 334152 149426 334332 149514
rect 334440 149426 334620 149514
rect 334728 149426 334908 149514
rect 335016 149426 335196 149514
rect 335304 149426 335484 149514
rect 335592 149426 335772 149514
rect 335880 149426 336060 149514
rect 336314 149426 336494 149514
rect 336602 149426 336782 149514
rect 336890 149426 337070 149514
rect 337178 149426 337358 149514
rect 337466 149426 337646 149514
rect 337754 149426 337934 149514
rect 338042 149426 338222 149514
rect 338330 149426 338510 149514
rect 338764 149426 338944 149514
rect 339052 149426 339232 149514
rect 339340 149426 339520 149514
rect 339628 149426 339808 149514
rect 339916 149426 340096 149514
rect 340204 149426 340384 149514
rect 340492 149426 340672 149514
rect 340780 149426 340960 149514
rect 341214 149426 341394 149514
rect 341502 149426 341682 149514
rect 341790 149426 341970 149514
rect 342078 149426 342258 149514
rect 342366 149426 342546 149514
rect 342654 149426 342834 149514
rect 342942 149426 343122 149514
rect 343230 149426 343410 149514
rect 343664 149426 343844 149514
rect 343952 149426 344132 149514
rect 344240 149426 344420 149514
rect 344528 149426 344708 149514
rect 344816 149426 344996 149514
rect 345104 149426 345284 149514
rect 345392 149426 345572 149514
rect 345680 149426 345860 149514
rect 346114 149426 346294 149514
rect 346402 149426 346582 149514
rect 346690 149426 346870 149514
rect 346978 149426 347158 149514
rect 347266 149426 347446 149514
rect 347554 149426 347734 149514
rect 347842 149426 348022 149514
rect 348130 149426 348310 149514
rect 348564 149426 348744 149514
rect 348852 149426 349032 149514
rect 349140 149426 349320 149514
rect 349428 149426 349608 149514
rect 349716 149426 349896 149514
rect 350004 149426 350184 149514
rect 350292 149426 350472 149514
rect 350580 149426 350760 149514
rect 351014 149426 351194 149514
rect 351302 149426 351482 149514
rect 351590 149426 351770 149514
rect 351878 149426 352058 149514
rect 352166 149426 352346 149514
rect 352454 149426 352634 149514
rect 352742 149426 352922 149514
rect 353030 149426 353210 149514
rect 353464 149426 353644 149514
rect 353752 149426 353932 149514
rect 354040 149426 354220 149514
rect 354328 149426 354508 149514
rect 354616 149426 354796 149514
rect 354904 149426 355084 149514
rect 355192 149426 355372 149514
rect 355480 149426 355660 149514
rect 355914 149426 356094 149514
rect 356202 149426 356382 149514
rect 356490 149426 356670 149514
rect 356778 149426 356958 149514
rect 357066 149426 357246 149514
rect 357354 149426 357534 149514
rect 357642 149426 357822 149514
rect 357930 149426 358110 149514
rect 358364 149426 358544 149514
rect 358652 149426 358832 149514
rect 358940 149426 359120 149514
rect 359228 149426 359408 149514
rect 359516 149426 359696 149514
rect 359804 149426 359984 149514
rect 360092 149426 360272 149514
rect 360380 149426 360560 149514
rect 360814 149426 360994 149514
rect 361102 149426 361282 149514
rect 361390 149426 361570 149514
rect 361678 149426 361858 149514
rect 361966 149426 362146 149514
rect 362254 149426 362434 149514
rect 362542 149426 362722 149514
rect 362830 149426 363010 149514
rect 363264 149426 363444 149514
rect 363552 149426 363732 149514
rect 363840 149426 364020 149514
rect 364128 149426 364308 149514
rect 364416 149426 364596 149514
rect 364704 149426 364884 149514
rect 364992 149426 365172 149514
rect 365280 149426 365460 149514
rect 365714 149426 365894 149514
rect 366002 149426 366182 149514
rect 366290 149426 366470 149514
rect 366578 149426 366758 149514
rect 366866 149426 367046 149514
rect 367154 149426 367334 149514
rect 367442 149426 367622 149514
rect 367730 149426 367910 149514
rect 243214 148950 243394 149038
rect 243502 148950 243682 149038
rect 243790 148950 243970 149038
rect 244078 148950 244258 149038
rect 244366 148950 244546 149038
rect 244654 148950 244834 149038
rect 244942 148950 245122 149038
rect 245230 148950 245410 149038
rect 245664 148950 245844 149038
rect 245952 148950 246132 149038
rect 246240 148950 246420 149038
rect 246528 148950 246708 149038
rect 246816 148950 246996 149038
rect 247104 148950 247284 149038
rect 247392 148950 247572 149038
rect 247680 148950 247860 149038
rect 248114 148950 248294 149038
rect 248402 148950 248582 149038
rect 248690 148950 248870 149038
rect 248978 148950 249158 149038
rect 249266 148950 249446 149038
rect 249554 148950 249734 149038
rect 249842 148950 250022 149038
rect 250130 148950 250310 149038
rect 250564 148950 250744 149038
rect 250852 148950 251032 149038
rect 251140 148950 251320 149038
rect 251428 148950 251608 149038
rect 251716 148950 251896 149038
rect 252004 148950 252184 149038
rect 252292 148950 252472 149038
rect 252580 148950 252760 149038
rect 253014 148950 253194 149038
rect 253302 148950 253482 149038
rect 253590 148950 253770 149038
rect 253878 148950 254058 149038
rect 254166 148950 254346 149038
rect 254454 148950 254634 149038
rect 254742 148950 254922 149038
rect 255030 148950 255210 149038
rect 255464 148950 255644 149038
rect 255752 148950 255932 149038
rect 256040 148950 256220 149038
rect 256328 148950 256508 149038
rect 256616 148950 256796 149038
rect 256904 148950 257084 149038
rect 257192 148950 257372 149038
rect 257480 148950 257660 149038
rect 257914 148950 258094 149038
rect 258202 148950 258382 149038
rect 258490 148950 258670 149038
rect 258778 148950 258958 149038
rect 259066 148950 259246 149038
rect 259354 148950 259534 149038
rect 259642 148950 259822 149038
rect 259930 148950 260110 149038
rect 260364 148950 260544 149038
rect 260652 148950 260832 149038
rect 260940 148950 261120 149038
rect 261228 148950 261408 149038
rect 261516 148950 261696 149038
rect 261804 148950 261984 149038
rect 262092 148950 262272 149038
rect 262380 148950 262560 149038
rect 262814 148950 262994 149038
rect 263102 148950 263282 149038
rect 263390 148950 263570 149038
rect 263678 148950 263858 149038
rect 263966 148950 264146 149038
rect 264254 148950 264434 149038
rect 264542 148950 264722 149038
rect 264830 148950 265010 149038
rect 265264 148950 265444 149038
rect 265552 148950 265732 149038
rect 265840 148950 266020 149038
rect 266128 148950 266308 149038
rect 266416 148950 266596 149038
rect 266704 148950 266884 149038
rect 266992 148950 267172 149038
rect 267280 148950 267460 149038
rect 267714 148950 267894 149038
rect 268002 148950 268182 149038
rect 268290 148950 268470 149038
rect 268578 148950 268758 149038
rect 268866 148950 269046 149038
rect 269154 148950 269334 149038
rect 269442 148950 269622 149038
rect 269730 148950 269910 149038
rect 270164 148950 270344 149038
rect 270452 148950 270632 149038
rect 270740 148950 270920 149038
rect 271028 148950 271208 149038
rect 271316 148950 271496 149038
rect 271604 148950 271784 149038
rect 271892 148950 272072 149038
rect 272180 148950 272360 149038
rect 272614 148950 272794 149038
rect 272902 148950 273082 149038
rect 273190 148950 273370 149038
rect 273478 148950 273658 149038
rect 273766 148950 273946 149038
rect 274054 148950 274234 149038
rect 274342 148950 274522 149038
rect 274630 148950 274810 149038
rect 275064 148950 275244 149038
rect 275352 148950 275532 149038
rect 275640 148950 275820 149038
rect 275928 148950 276108 149038
rect 276216 148950 276396 149038
rect 276504 148950 276684 149038
rect 276792 148950 276972 149038
rect 277080 148950 277260 149038
rect 277514 148950 277694 149038
rect 277802 148950 277982 149038
rect 278090 148950 278270 149038
rect 278378 148950 278558 149038
rect 278666 148950 278846 149038
rect 278954 148950 279134 149038
rect 279242 148950 279422 149038
rect 279530 148950 279710 149038
rect 279964 148950 280144 149038
rect 280252 148950 280432 149038
rect 280540 148950 280720 149038
rect 280828 148950 281008 149038
rect 281116 148950 281296 149038
rect 281404 148950 281584 149038
rect 281692 148950 281872 149038
rect 281980 148950 282160 149038
rect 282414 148950 282594 149038
rect 282702 148950 282882 149038
rect 282990 148950 283170 149038
rect 283278 148950 283458 149038
rect 283566 148950 283746 149038
rect 283854 148950 284034 149038
rect 284142 148950 284322 149038
rect 284430 148950 284610 149038
rect 284864 148950 285044 149038
rect 285152 148950 285332 149038
rect 285440 148950 285620 149038
rect 285728 148950 285908 149038
rect 286016 148950 286196 149038
rect 286304 148950 286484 149038
rect 286592 148950 286772 149038
rect 286880 148950 287060 149038
rect 287314 148950 287494 149038
rect 287602 148950 287782 149038
rect 287890 148950 288070 149038
rect 288178 148950 288358 149038
rect 288466 148950 288646 149038
rect 288754 148950 288934 149038
rect 289042 148950 289222 149038
rect 289330 148950 289510 149038
rect 289764 148950 289944 149038
rect 290052 148950 290232 149038
rect 290340 148950 290520 149038
rect 290628 148950 290808 149038
rect 290916 148950 291096 149038
rect 291204 148950 291384 149038
rect 291492 148950 291672 149038
rect 291780 148950 291960 149038
rect 292214 148950 292394 149038
rect 292502 148950 292682 149038
rect 292790 148950 292970 149038
rect 293078 148950 293258 149038
rect 293366 148950 293546 149038
rect 293654 148950 293834 149038
rect 293942 148950 294122 149038
rect 294230 148950 294410 149038
rect 294664 148950 294844 149038
rect 294952 148950 295132 149038
rect 295240 148950 295420 149038
rect 295528 148950 295708 149038
rect 295816 148950 295996 149038
rect 296104 148950 296284 149038
rect 296392 148950 296572 149038
rect 296680 148950 296860 149038
rect 297114 148950 297294 149038
rect 297402 148950 297582 149038
rect 297690 148950 297870 149038
rect 297978 148950 298158 149038
rect 298266 148950 298446 149038
rect 298554 148950 298734 149038
rect 298842 148950 299022 149038
rect 299130 148950 299310 149038
rect 299564 148950 299744 149038
rect 299852 148950 300032 149038
rect 300140 148950 300320 149038
rect 300428 148950 300608 149038
rect 300716 148950 300896 149038
rect 301004 148950 301184 149038
rect 301292 148950 301472 149038
rect 301580 148950 301760 149038
rect 302014 148950 302194 149038
rect 302302 148950 302482 149038
rect 302590 148950 302770 149038
rect 302878 148950 303058 149038
rect 303166 148950 303346 149038
rect 303454 148950 303634 149038
rect 303742 148950 303922 149038
rect 304030 148950 304210 149038
rect 304464 148950 304644 149038
rect 304752 148950 304932 149038
rect 305040 148950 305220 149038
rect 305328 148950 305508 149038
rect 305616 148950 305796 149038
rect 305904 148950 306084 149038
rect 306192 148950 306372 149038
rect 306480 148950 306660 149038
rect 306914 148950 307094 149038
rect 307202 148950 307382 149038
rect 307490 148950 307670 149038
rect 307778 148950 307958 149038
rect 308066 148950 308246 149038
rect 308354 148950 308534 149038
rect 308642 148950 308822 149038
rect 308930 148950 309110 149038
rect 309364 148950 309544 149038
rect 309652 148950 309832 149038
rect 309940 148950 310120 149038
rect 310228 148950 310408 149038
rect 310516 148950 310696 149038
rect 310804 148950 310984 149038
rect 311092 148950 311272 149038
rect 311380 148950 311560 149038
rect 311814 148950 311994 149038
rect 312102 148950 312282 149038
rect 312390 148950 312570 149038
rect 312678 148950 312858 149038
rect 312966 148950 313146 149038
rect 313254 148950 313434 149038
rect 313542 148950 313722 149038
rect 313830 148950 314010 149038
rect 314264 148950 314444 149038
rect 314552 148950 314732 149038
rect 314840 148950 315020 149038
rect 315128 148950 315308 149038
rect 315416 148950 315596 149038
rect 315704 148950 315884 149038
rect 315992 148950 316172 149038
rect 316280 148950 316460 149038
rect 316714 148950 316894 149038
rect 317002 148950 317182 149038
rect 317290 148950 317470 149038
rect 317578 148950 317758 149038
rect 317866 148950 318046 149038
rect 318154 148950 318334 149038
rect 318442 148950 318622 149038
rect 318730 148950 318910 149038
rect 319164 148950 319344 149038
rect 319452 148950 319632 149038
rect 319740 148950 319920 149038
rect 320028 148950 320208 149038
rect 320316 148950 320496 149038
rect 320604 148950 320784 149038
rect 320892 148950 321072 149038
rect 321180 148950 321360 149038
rect 321614 148950 321794 149038
rect 321902 148950 322082 149038
rect 322190 148950 322370 149038
rect 322478 148950 322658 149038
rect 322766 148950 322946 149038
rect 323054 148950 323234 149038
rect 323342 148950 323522 149038
rect 323630 148950 323810 149038
rect 324064 148950 324244 149038
rect 324352 148950 324532 149038
rect 324640 148950 324820 149038
rect 324928 148950 325108 149038
rect 325216 148950 325396 149038
rect 325504 148950 325684 149038
rect 325792 148950 325972 149038
rect 326080 148950 326260 149038
rect 326514 148950 326694 149038
rect 326802 148950 326982 149038
rect 327090 148950 327270 149038
rect 327378 148950 327558 149038
rect 327666 148950 327846 149038
rect 327954 148950 328134 149038
rect 328242 148950 328422 149038
rect 328530 148950 328710 149038
rect 328964 148950 329144 149038
rect 329252 148950 329432 149038
rect 329540 148950 329720 149038
rect 329828 148950 330008 149038
rect 330116 148950 330296 149038
rect 330404 148950 330584 149038
rect 330692 148950 330872 149038
rect 330980 148950 331160 149038
rect 331414 148950 331594 149038
rect 331702 148950 331882 149038
rect 331990 148950 332170 149038
rect 332278 148950 332458 149038
rect 332566 148950 332746 149038
rect 332854 148950 333034 149038
rect 333142 148950 333322 149038
rect 333430 148950 333610 149038
rect 333864 148950 334044 149038
rect 334152 148950 334332 149038
rect 334440 148950 334620 149038
rect 334728 148950 334908 149038
rect 335016 148950 335196 149038
rect 335304 148950 335484 149038
rect 335592 148950 335772 149038
rect 335880 148950 336060 149038
rect 336314 148950 336494 149038
rect 336602 148950 336782 149038
rect 336890 148950 337070 149038
rect 337178 148950 337358 149038
rect 337466 148950 337646 149038
rect 337754 148950 337934 149038
rect 338042 148950 338222 149038
rect 338330 148950 338510 149038
rect 338764 148950 338944 149038
rect 339052 148950 339232 149038
rect 339340 148950 339520 149038
rect 339628 148950 339808 149038
rect 339916 148950 340096 149038
rect 340204 148950 340384 149038
rect 340492 148950 340672 149038
rect 340780 148950 340960 149038
rect 341214 148950 341394 149038
rect 341502 148950 341682 149038
rect 341790 148950 341970 149038
rect 342078 148950 342258 149038
rect 342366 148950 342546 149038
rect 342654 148950 342834 149038
rect 342942 148950 343122 149038
rect 343230 148950 343410 149038
rect 343664 148950 343844 149038
rect 343952 148950 344132 149038
rect 344240 148950 344420 149038
rect 344528 148950 344708 149038
rect 344816 148950 344996 149038
rect 345104 148950 345284 149038
rect 345392 148950 345572 149038
rect 345680 148950 345860 149038
rect 346114 148950 346294 149038
rect 346402 148950 346582 149038
rect 346690 148950 346870 149038
rect 346978 148950 347158 149038
rect 347266 148950 347446 149038
rect 347554 148950 347734 149038
rect 347842 148950 348022 149038
rect 348130 148950 348310 149038
rect 348564 148950 348744 149038
rect 348852 148950 349032 149038
rect 349140 148950 349320 149038
rect 349428 148950 349608 149038
rect 349716 148950 349896 149038
rect 350004 148950 350184 149038
rect 350292 148950 350472 149038
rect 350580 148950 350760 149038
rect 351014 148950 351194 149038
rect 351302 148950 351482 149038
rect 351590 148950 351770 149038
rect 351878 148950 352058 149038
rect 352166 148950 352346 149038
rect 352454 148950 352634 149038
rect 352742 148950 352922 149038
rect 353030 148950 353210 149038
rect 353464 148950 353644 149038
rect 353752 148950 353932 149038
rect 354040 148950 354220 149038
rect 354328 148950 354508 149038
rect 354616 148950 354796 149038
rect 354904 148950 355084 149038
rect 355192 148950 355372 149038
rect 355480 148950 355660 149038
rect 355914 148950 356094 149038
rect 356202 148950 356382 149038
rect 356490 148950 356670 149038
rect 356778 148950 356958 149038
rect 357066 148950 357246 149038
rect 357354 148950 357534 149038
rect 357642 148950 357822 149038
rect 357930 148950 358110 149038
rect 358364 148950 358544 149038
rect 358652 148950 358832 149038
rect 358940 148950 359120 149038
rect 359228 148950 359408 149038
rect 359516 148950 359696 149038
rect 359804 148950 359984 149038
rect 360092 148950 360272 149038
rect 360380 148950 360560 149038
rect 360814 148950 360994 149038
rect 361102 148950 361282 149038
rect 361390 148950 361570 149038
rect 361678 148950 361858 149038
rect 361966 148950 362146 149038
rect 362254 148950 362434 149038
rect 362542 148950 362722 149038
rect 362830 148950 363010 149038
rect 363264 148950 363444 149038
rect 363552 148950 363732 149038
rect 363840 148950 364020 149038
rect 364128 148950 364308 149038
rect 364416 148950 364596 149038
rect 364704 148950 364884 149038
rect 364992 148950 365172 149038
rect 365280 148950 365460 149038
rect 365714 148950 365894 149038
rect 366002 148950 366182 149038
rect 366290 148950 366470 149038
rect 366578 148950 366758 149038
rect 366866 148950 367046 149038
rect 367154 148950 367334 149038
rect 367442 148950 367622 149038
rect 367730 148950 367910 149038
rect 243214 148476 243394 148564
rect 243502 148476 243682 148564
rect 243790 148476 243970 148564
rect 244078 148476 244258 148564
rect 244366 148476 244546 148564
rect 244654 148476 244834 148564
rect 244942 148476 245122 148564
rect 245230 148476 245410 148564
rect 245664 148476 245844 148564
rect 245952 148476 246132 148564
rect 246240 148476 246420 148564
rect 246528 148476 246708 148564
rect 246816 148476 246996 148564
rect 247104 148476 247284 148564
rect 247392 148476 247572 148564
rect 247680 148476 247860 148564
rect 248114 148476 248294 148564
rect 248402 148476 248582 148564
rect 248690 148476 248870 148564
rect 248978 148476 249158 148564
rect 249266 148476 249446 148564
rect 249554 148476 249734 148564
rect 249842 148476 250022 148564
rect 250130 148476 250310 148564
rect 250564 148476 250744 148564
rect 250852 148476 251032 148564
rect 251140 148476 251320 148564
rect 251428 148476 251608 148564
rect 251716 148476 251896 148564
rect 252004 148476 252184 148564
rect 252292 148476 252472 148564
rect 252580 148476 252760 148564
rect 253014 148476 253194 148564
rect 253302 148476 253482 148564
rect 253590 148476 253770 148564
rect 253878 148476 254058 148564
rect 254166 148476 254346 148564
rect 254454 148476 254634 148564
rect 254742 148476 254922 148564
rect 255030 148476 255210 148564
rect 255464 148476 255644 148564
rect 255752 148476 255932 148564
rect 256040 148476 256220 148564
rect 256328 148476 256508 148564
rect 256616 148476 256796 148564
rect 256904 148476 257084 148564
rect 257192 148476 257372 148564
rect 257480 148476 257660 148564
rect 257914 148476 258094 148564
rect 258202 148476 258382 148564
rect 258490 148476 258670 148564
rect 258778 148476 258958 148564
rect 259066 148476 259246 148564
rect 259354 148476 259534 148564
rect 259642 148476 259822 148564
rect 259930 148476 260110 148564
rect 260364 148476 260544 148564
rect 260652 148476 260832 148564
rect 260940 148476 261120 148564
rect 261228 148476 261408 148564
rect 261516 148476 261696 148564
rect 261804 148476 261984 148564
rect 262092 148476 262272 148564
rect 262380 148476 262560 148564
rect 262814 148476 262994 148564
rect 263102 148476 263282 148564
rect 263390 148476 263570 148564
rect 263678 148476 263858 148564
rect 263966 148476 264146 148564
rect 264254 148476 264434 148564
rect 264542 148476 264722 148564
rect 264830 148476 265010 148564
rect 265264 148476 265444 148564
rect 265552 148476 265732 148564
rect 265840 148476 266020 148564
rect 266128 148476 266308 148564
rect 266416 148476 266596 148564
rect 266704 148476 266884 148564
rect 266992 148476 267172 148564
rect 267280 148476 267460 148564
rect 267714 148476 267894 148564
rect 268002 148476 268182 148564
rect 268290 148476 268470 148564
rect 268578 148476 268758 148564
rect 268866 148476 269046 148564
rect 269154 148476 269334 148564
rect 269442 148476 269622 148564
rect 269730 148476 269910 148564
rect 270164 148476 270344 148564
rect 270452 148476 270632 148564
rect 270740 148476 270920 148564
rect 271028 148476 271208 148564
rect 271316 148476 271496 148564
rect 271604 148476 271784 148564
rect 271892 148476 272072 148564
rect 272180 148476 272360 148564
rect 272614 148476 272794 148564
rect 272902 148476 273082 148564
rect 273190 148476 273370 148564
rect 273478 148476 273658 148564
rect 273766 148476 273946 148564
rect 274054 148476 274234 148564
rect 274342 148476 274522 148564
rect 274630 148476 274810 148564
rect 275064 148476 275244 148564
rect 275352 148476 275532 148564
rect 275640 148476 275820 148564
rect 275928 148476 276108 148564
rect 276216 148476 276396 148564
rect 276504 148476 276684 148564
rect 276792 148476 276972 148564
rect 277080 148476 277260 148564
rect 277514 148476 277694 148564
rect 277802 148476 277982 148564
rect 278090 148476 278270 148564
rect 278378 148476 278558 148564
rect 278666 148476 278846 148564
rect 278954 148476 279134 148564
rect 279242 148476 279422 148564
rect 279530 148476 279710 148564
rect 279964 148476 280144 148564
rect 280252 148476 280432 148564
rect 280540 148476 280720 148564
rect 280828 148476 281008 148564
rect 281116 148476 281296 148564
rect 281404 148476 281584 148564
rect 281692 148476 281872 148564
rect 281980 148476 282160 148564
rect 282414 148476 282594 148564
rect 282702 148476 282882 148564
rect 282990 148476 283170 148564
rect 283278 148476 283458 148564
rect 283566 148476 283746 148564
rect 283854 148476 284034 148564
rect 284142 148476 284322 148564
rect 284430 148476 284610 148564
rect 284864 148476 285044 148564
rect 285152 148476 285332 148564
rect 285440 148476 285620 148564
rect 285728 148476 285908 148564
rect 286016 148476 286196 148564
rect 286304 148476 286484 148564
rect 286592 148476 286772 148564
rect 286880 148476 287060 148564
rect 287314 148476 287494 148564
rect 287602 148476 287782 148564
rect 287890 148476 288070 148564
rect 288178 148476 288358 148564
rect 288466 148476 288646 148564
rect 288754 148476 288934 148564
rect 289042 148476 289222 148564
rect 289330 148476 289510 148564
rect 289764 148476 289944 148564
rect 290052 148476 290232 148564
rect 290340 148476 290520 148564
rect 290628 148476 290808 148564
rect 290916 148476 291096 148564
rect 291204 148476 291384 148564
rect 291492 148476 291672 148564
rect 291780 148476 291960 148564
rect 292214 148476 292394 148564
rect 292502 148476 292682 148564
rect 292790 148476 292970 148564
rect 293078 148476 293258 148564
rect 293366 148476 293546 148564
rect 293654 148476 293834 148564
rect 293942 148476 294122 148564
rect 294230 148476 294410 148564
rect 294664 148476 294844 148564
rect 294952 148476 295132 148564
rect 295240 148476 295420 148564
rect 295528 148476 295708 148564
rect 295816 148476 295996 148564
rect 296104 148476 296284 148564
rect 296392 148476 296572 148564
rect 296680 148476 296860 148564
rect 297114 148476 297294 148564
rect 297402 148476 297582 148564
rect 297690 148476 297870 148564
rect 297978 148476 298158 148564
rect 298266 148476 298446 148564
rect 298554 148476 298734 148564
rect 298842 148476 299022 148564
rect 299130 148476 299310 148564
rect 299564 148476 299744 148564
rect 299852 148476 300032 148564
rect 300140 148476 300320 148564
rect 300428 148476 300608 148564
rect 300716 148476 300896 148564
rect 301004 148476 301184 148564
rect 301292 148476 301472 148564
rect 301580 148476 301760 148564
rect 302014 148476 302194 148564
rect 302302 148476 302482 148564
rect 302590 148476 302770 148564
rect 302878 148476 303058 148564
rect 303166 148476 303346 148564
rect 303454 148476 303634 148564
rect 303742 148476 303922 148564
rect 304030 148476 304210 148564
rect 304464 148476 304644 148564
rect 304752 148476 304932 148564
rect 305040 148476 305220 148564
rect 305328 148476 305508 148564
rect 305616 148476 305796 148564
rect 305904 148476 306084 148564
rect 306192 148476 306372 148564
rect 306480 148476 306660 148564
rect 306914 148476 307094 148564
rect 307202 148476 307382 148564
rect 307490 148476 307670 148564
rect 307778 148476 307958 148564
rect 308066 148476 308246 148564
rect 308354 148476 308534 148564
rect 308642 148476 308822 148564
rect 308930 148476 309110 148564
rect 309364 148476 309544 148564
rect 309652 148476 309832 148564
rect 309940 148476 310120 148564
rect 310228 148476 310408 148564
rect 310516 148476 310696 148564
rect 310804 148476 310984 148564
rect 311092 148476 311272 148564
rect 311380 148476 311560 148564
rect 311814 148476 311994 148564
rect 312102 148476 312282 148564
rect 312390 148476 312570 148564
rect 312678 148476 312858 148564
rect 312966 148476 313146 148564
rect 313254 148476 313434 148564
rect 313542 148476 313722 148564
rect 313830 148476 314010 148564
rect 314264 148476 314444 148564
rect 314552 148476 314732 148564
rect 314840 148476 315020 148564
rect 315128 148476 315308 148564
rect 315416 148476 315596 148564
rect 315704 148476 315884 148564
rect 315992 148476 316172 148564
rect 316280 148476 316460 148564
rect 316714 148476 316894 148564
rect 317002 148476 317182 148564
rect 317290 148476 317470 148564
rect 317578 148476 317758 148564
rect 317866 148476 318046 148564
rect 318154 148476 318334 148564
rect 318442 148476 318622 148564
rect 318730 148476 318910 148564
rect 319164 148476 319344 148564
rect 319452 148476 319632 148564
rect 319740 148476 319920 148564
rect 320028 148476 320208 148564
rect 320316 148476 320496 148564
rect 320604 148476 320784 148564
rect 320892 148476 321072 148564
rect 321180 148476 321360 148564
rect 321614 148476 321794 148564
rect 321902 148476 322082 148564
rect 322190 148476 322370 148564
rect 322478 148476 322658 148564
rect 322766 148476 322946 148564
rect 323054 148476 323234 148564
rect 323342 148476 323522 148564
rect 323630 148476 323810 148564
rect 324064 148476 324244 148564
rect 324352 148476 324532 148564
rect 324640 148476 324820 148564
rect 324928 148476 325108 148564
rect 325216 148476 325396 148564
rect 325504 148476 325684 148564
rect 325792 148476 325972 148564
rect 326080 148476 326260 148564
rect 326514 148476 326694 148564
rect 326802 148476 326982 148564
rect 327090 148476 327270 148564
rect 327378 148476 327558 148564
rect 327666 148476 327846 148564
rect 327954 148476 328134 148564
rect 328242 148476 328422 148564
rect 328530 148476 328710 148564
rect 328964 148476 329144 148564
rect 329252 148476 329432 148564
rect 329540 148476 329720 148564
rect 329828 148476 330008 148564
rect 330116 148476 330296 148564
rect 330404 148476 330584 148564
rect 330692 148476 330872 148564
rect 330980 148476 331160 148564
rect 331414 148476 331594 148564
rect 331702 148476 331882 148564
rect 331990 148476 332170 148564
rect 332278 148476 332458 148564
rect 332566 148476 332746 148564
rect 332854 148476 333034 148564
rect 333142 148476 333322 148564
rect 333430 148476 333610 148564
rect 333864 148476 334044 148564
rect 334152 148476 334332 148564
rect 334440 148476 334620 148564
rect 334728 148476 334908 148564
rect 335016 148476 335196 148564
rect 335304 148476 335484 148564
rect 335592 148476 335772 148564
rect 335880 148476 336060 148564
rect 336314 148476 336494 148564
rect 336602 148476 336782 148564
rect 336890 148476 337070 148564
rect 337178 148476 337358 148564
rect 337466 148476 337646 148564
rect 337754 148476 337934 148564
rect 338042 148476 338222 148564
rect 338330 148476 338510 148564
rect 338764 148476 338944 148564
rect 339052 148476 339232 148564
rect 339340 148476 339520 148564
rect 339628 148476 339808 148564
rect 339916 148476 340096 148564
rect 340204 148476 340384 148564
rect 340492 148476 340672 148564
rect 340780 148476 340960 148564
rect 341214 148476 341394 148564
rect 341502 148476 341682 148564
rect 341790 148476 341970 148564
rect 342078 148476 342258 148564
rect 342366 148476 342546 148564
rect 342654 148476 342834 148564
rect 342942 148476 343122 148564
rect 343230 148476 343410 148564
rect 343664 148476 343844 148564
rect 343952 148476 344132 148564
rect 344240 148476 344420 148564
rect 344528 148476 344708 148564
rect 344816 148476 344996 148564
rect 345104 148476 345284 148564
rect 345392 148476 345572 148564
rect 345680 148476 345860 148564
rect 346114 148476 346294 148564
rect 346402 148476 346582 148564
rect 346690 148476 346870 148564
rect 346978 148476 347158 148564
rect 347266 148476 347446 148564
rect 347554 148476 347734 148564
rect 347842 148476 348022 148564
rect 348130 148476 348310 148564
rect 348564 148476 348744 148564
rect 348852 148476 349032 148564
rect 349140 148476 349320 148564
rect 349428 148476 349608 148564
rect 349716 148476 349896 148564
rect 350004 148476 350184 148564
rect 350292 148476 350472 148564
rect 350580 148476 350760 148564
rect 351014 148476 351194 148564
rect 351302 148476 351482 148564
rect 351590 148476 351770 148564
rect 351878 148476 352058 148564
rect 352166 148476 352346 148564
rect 352454 148476 352634 148564
rect 352742 148476 352922 148564
rect 353030 148476 353210 148564
rect 353464 148476 353644 148564
rect 353752 148476 353932 148564
rect 354040 148476 354220 148564
rect 354328 148476 354508 148564
rect 354616 148476 354796 148564
rect 354904 148476 355084 148564
rect 355192 148476 355372 148564
rect 355480 148476 355660 148564
rect 355914 148476 356094 148564
rect 356202 148476 356382 148564
rect 356490 148476 356670 148564
rect 356778 148476 356958 148564
rect 357066 148476 357246 148564
rect 357354 148476 357534 148564
rect 357642 148476 357822 148564
rect 357930 148476 358110 148564
rect 358364 148476 358544 148564
rect 358652 148476 358832 148564
rect 358940 148476 359120 148564
rect 359228 148476 359408 148564
rect 359516 148476 359696 148564
rect 359804 148476 359984 148564
rect 360092 148476 360272 148564
rect 360380 148476 360560 148564
rect 360814 148476 360994 148564
rect 361102 148476 361282 148564
rect 361390 148476 361570 148564
rect 361678 148476 361858 148564
rect 361966 148476 362146 148564
rect 362254 148476 362434 148564
rect 362542 148476 362722 148564
rect 362830 148476 363010 148564
rect 363264 148476 363444 148564
rect 363552 148476 363732 148564
rect 363840 148476 364020 148564
rect 364128 148476 364308 148564
rect 364416 148476 364596 148564
rect 364704 148476 364884 148564
rect 364992 148476 365172 148564
rect 365280 148476 365460 148564
rect 365714 148476 365894 148564
rect 366002 148476 366182 148564
rect 366290 148476 366470 148564
rect 366578 148476 366758 148564
rect 366866 148476 367046 148564
rect 367154 148476 367334 148564
rect 367442 148476 367622 148564
rect 367730 148476 367910 148564
rect 243214 148000 243394 148088
rect 243502 148000 243682 148088
rect 243790 148000 243970 148088
rect 244078 148000 244258 148088
rect 244366 148000 244546 148088
rect 244654 148000 244834 148088
rect 244942 148000 245122 148088
rect 245230 148000 245410 148088
rect 245664 148000 245844 148088
rect 245952 148000 246132 148088
rect 246240 148000 246420 148088
rect 246528 148000 246708 148088
rect 246816 148000 246996 148088
rect 247104 148000 247284 148088
rect 247392 148000 247572 148088
rect 247680 148000 247860 148088
rect 248114 148000 248294 148088
rect 248402 148000 248582 148088
rect 248690 148000 248870 148088
rect 248978 148000 249158 148088
rect 249266 148000 249446 148088
rect 249554 148000 249734 148088
rect 249842 148000 250022 148088
rect 250130 148000 250310 148088
rect 250564 148000 250744 148088
rect 250852 148000 251032 148088
rect 251140 148000 251320 148088
rect 251428 148000 251608 148088
rect 251716 148000 251896 148088
rect 252004 148000 252184 148088
rect 252292 148000 252472 148088
rect 252580 148000 252760 148088
rect 253014 148000 253194 148088
rect 253302 148000 253482 148088
rect 253590 148000 253770 148088
rect 253878 148000 254058 148088
rect 254166 148000 254346 148088
rect 254454 148000 254634 148088
rect 254742 148000 254922 148088
rect 255030 148000 255210 148088
rect 255464 148000 255644 148088
rect 255752 148000 255932 148088
rect 256040 148000 256220 148088
rect 256328 148000 256508 148088
rect 256616 148000 256796 148088
rect 256904 148000 257084 148088
rect 257192 148000 257372 148088
rect 257480 148000 257660 148088
rect 257914 148000 258094 148088
rect 258202 148000 258382 148088
rect 258490 148000 258670 148088
rect 258778 148000 258958 148088
rect 259066 148000 259246 148088
rect 259354 148000 259534 148088
rect 259642 148000 259822 148088
rect 259930 148000 260110 148088
rect 260364 148000 260544 148088
rect 260652 148000 260832 148088
rect 260940 148000 261120 148088
rect 261228 148000 261408 148088
rect 261516 148000 261696 148088
rect 261804 148000 261984 148088
rect 262092 148000 262272 148088
rect 262380 148000 262560 148088
rect 262814 148000 262994 148088
rect 263102 148000 263282 148088
rect 263390 148000 263570 148088
rect 263678 148000 263858 148088
rect 263966 148000 264146 148088
rect 264254 148000 264434 148088
rect 264542 148000 264722 148088
rect 264830 148000 265010 148088
rect 265264 148000 265444 148088
rect 265552 148000 265732 148088
rect 265840 148000 266020 148088
rect 266128 148000 266308 148088
rect 266416 148000 266596 148088
rect 266704 148000 266884 148088
rect 266992 148000 267172 148088
rect 267280 148000 267460 148088
rect 267714 148000 267894 148088
rect 268002 148000 268182 148088
rect 268290 148000 268470 148088
rect 268578 148000 268758 148088
rect 268866 148000 269046 148088
rect 269154 148000 269334 148088
rect 269442 148000 269622 148088
rect 269730 148000 269910 148088
rect 270164 148000 270344 148088
rect 270452 148000 270632 148088
rect 270740 148000 270920 148088
rect 271028 148000 271208 148088
rect 271316 148000 271496 148088
rect 271604 148000 271784 148088
rect 271892 148000 272072 148088
rect 272180 148000 272360 148088
rect 272614 148000 272794 148088
rect 272902 148000 273082 148088
rect 273190 148000 273370 148088
rect 273478 148000 273658 148088
rect 273766 148000 273946 148088
rect 274054 148000 274234 148088
rect 274342 148000 274522 148088
rect 274630 148000 274810 148088
rect 275064 148000 275244 148088
rect 275352 148000 275532 148088
rect 275640 148000 275820 148088
rect 275928 148000 276108 148088
rect 276216 148000 276396 148088
rect 276504 148000 276684 148088
rect 276792 148000 276972 148088
rect 277080 148000 277260 148088
rect 277514 148000 277694 148088
rect 277802 148000 277982 148088
rect 278090 148000 278270 148088
rect 278378 148000 278558 148088
rect 278666 148000 278846 148088
rect 278954 148000 279134 148088
rect 279242 148000 279422 148088
rect 279530 148000 279710 148088
rect 279964 148000 280144 148088
rect 280252 148000 280432 148088
rect 280540 148000 280720 148088
rect 280828 148000 281008 148088
rect 281116 148000 281296 148088
rect 281404 148000 281584 148088
rect 281692 148000 281872 148088
rect 281980 148000 282160 148088
rect 282414 148000 282594 148088
rect 282702 148000 282882 148088
rect 282990 148000 283170 148088
rect 283278 148000 283458 148088
rect 283566 148000 283746 148088
rect 283854 148000 284034 148088
rect 284142 148000 284322 148088
rect 284430 148000 284610 148088
rect 284864 148000 285044 148088
rect 285152 148000 285332 148088
rect 285440 148000 285620 148088
rect 285728 148000 285908 148088
rect 286016 148000 286196 148088
rect 286304 148000 286484 148088
rect 286592 148000 286772 148088
rect 286880 148000 287060 148088
rect 287314 148000 287494 148088
rect 287602 148000 287782 148088
rect 287890 148000 288070 148088
rect 288178 148000 288358 148088
rect 288466 148000 288646 148088
rect 288754 148000 288934 148088
rect 289042 148000 289222 148088
rect 289330 148000 289510 148088
rect 289764 148000 289944 148088
rect 290052 148000 290232 148088
rect 290340 148000 290520 148088
rect 290628 148000 290808 148088
rect 290916 148000 291096 148088
rect 291204 148000 291384 148088
rect 291492 148000 291672 148088
rect 291780 148000 291960 148088
rect 292214 148000 292394 148088
rect 292502 148000 292682 148088
rect 292790 148000 292970 148088
rect 293078 148000 293258 148088
rect 293366 148000 293546 148088
rect 293654 148000 293834 148088
rect 293942 148000 294122 148088
rect 294230 148000 294410 148088
rect 294664 148000 294844 148088
rect 294952 148000 295132 148088
rect 295240 148000 295420 148088
rect 295528 148000 295708 148088
rect 295816 148000 295996 148088
rect 296104 148000 296284 148088
rect 296392 148000 296572 148088
rect 296680 148000 296860 148088
rect 297114 148000 297294 148088
rect 297402 148000 297582 148088
rect 297690 148000 297870 148088
rect 297978 148000 298158 148088
rect 298266 148000 298446 148088
rect 298554 148000 298734 148088
rect 298842 148000 299022 148088
rect 299130 148000 299310 148088
rect 299564 148000 299744 148088
rect 299852 148000 300032 148088
rect 300140 148000 300320 148088
rect 300428 148000 300608 148088
rect 300716 148000 300896 148088
rect 301004 148000 301184 148088
rect 301292 148000 301472 148088
rect 301580 148000 301760 148088
rect 302014 148000 302194 148088
rect 302302 148000 302482 148088
rect 302590 148000 302770 148088
rect 302878 148000 303058 148088
rect 303166 148000 303346 148088
rect 303454 148000 303634 148088
rect 303742 148000 303922 148088
rect 304030 148000 304210 148088
rect 304464 148000 304644 148088
rect 304752 148000 304932 148088
rect 305040 148000 305220 148088
rect 305328 148000 305508 148088
rect 305616 148000 305796 148088
rect 305904 148000 306084 148088
rect 306192 148000 306372 148088
rect 306480 148000 306660 148088
rect 306914 148000 307094 148088
rect 307202 148000 307382 148088
rect 307490 148000 307670 148088
rect 307778 148000 307958 148088
rect 308066 148000 308246 148088
rect 308354 148000 308534 148088
rect 308642 148000 308822 148088
rect 308930 148000 309110 148088
rect 309364 148000 309544 148088
rect 309652 148000 309832 148088
rect 309940 148000 310120 148088
rect 310228 148000 310408 148088
rect 310516 148000 310696 148088
rect 310804 148000 310984 148088
rect 311092 148000 311272 148088
rect 311380 148000 311560 148088
rect 311814 148000 311994 148088
rect 312102 148000 312282 148088
rect 312390 148000 312570 148088
rect 312678 148000 312858 148088
rect 312966 148000 313146 148088
rect 313254 148000 313434 148088
rect 313542 148000 313722 148088
rect 313830 148000 314010 148088
rect 314264 148000 314444 148088
rect 314552 148000 314732 148088
rect 314840 148000 315020 148088
rect 315128 148000 315308 148088
rect 315416 148000 315596 148088
rect 315704 148000 315884 148088
rect 315992 148000 316172 148088
rect 316280 148000 316460 148088
rect 316714 148000 316894 148088
rect 317002 148000 317182 148088
rect 317290 148000 317470 148088
rect 317578 148000 317758 148088
rect 317866 148000 318046 148088
rect 318154 148000 318334 148088
rect 318442 148000 318622 148088
rect 318730 148000 318910 148088
rect 319164 148000 319344 148088
rect 319452 148000 319632 148088
rect 319740 148000 319920 148088
rect 320028 148000 320208 148088
rect 320316 148000 320496 148088
rect 320604 148000 320784 148088
rect 320892 148000 321072 148088
rect 321180 148000 321360 148088
rect 321614 148000 321794 148088
rect 321902 148000 322082 148088
rect 322190 148000 322370 148088
rect 322478 148000 322658 148088
rect 322766 148000 322946 148088
rect 323054 148000 323234 148088
rect 323342 148000 323522 148088
rect 323630 148000 323810 148088
rect 324064 148000 324244 148088
rect 324352 148000 324532 148088
rect 324640 148000 324820 148088
rect 324928 148000 325108 148088
rect 325216 148000 325396 148088
rect 325504 148000 325684 148088
rect 325792 148000 325972 148088
rect 326080 148000 326260 148088
rect 326514 148000 326694 148088
rect 326802 148000 326982 148088
rect 327090 148000 327270 148088
rect 327378 148000 327558 148088
rect 327666 148000 327846 148088
rect 327954 148000 328134 148088
rect 328242 148000 328422 148088
rect 328530 148000 328710 148088
rect 328964 148000 329144 148088
rect 329252 148000 329432 148088
rect 329540 148000 329720 148088
rect 329828 148000 330008 148088
rect 330116 148000 330296 148088
rect 330404 148000 330584 148088
rect 330692 148000 330872 148088
rect 330980 148000 331160 148088
rect 331414 148000 331594 148088
rect 331702 148000 331882 148088
rect 331990 148000 332170 148088
rect 332278 148000 332458 148088
rect 332566 148000 332746 148088
rect 332854 148000 333034 148088
rect 333142 148000 333322 148088
rect 333430 148000 333610 148088
rect 333864 148000 334044 148088
rect 334152 148000 334332 148088
rect 334440 148000 334620 148088
rect 334728 148000 334908 148088
rect 335016 148000 335196 148088
rect 335304 148000 335484 148088
rect 335592 148000 335772 148088
rect 335880 148000 336060 148088
rect 336314 148000 336494 148088
rect 336602 148000 336782 148088
rect 336890 148000 337070 148088
rect 337178 148000 337358 148088
rect 337466 148000 337646 148088
rect 337754 148000 337934 148088
rect 338042 148000 338222 148088
rect 338330 148000 338510 148088
rect 338764 148000 338944 148088
rect 339052 148000 339232 148088
rect 339340 148000 339520 148088
rect 339628 148000 339808 148088
rect 339916 148000 340096 148088
rect 340204 148000 340384 148088
rect 340492 148000 340672 148088
rect 340780 148000 340960 148088
rect 341214 148000 341394 148088
rect 341502 148000 341682 148088
rect 341790 148000 341970 148088
rect 342078 148000 342258 148088
rect 342366 148000 342546 148088
rect 342654 148000 342834 148088
rect 342942 148000 343122 148088
rect 343230 148000 343410 148088
rect 343664 148000 343844 148088
rect 343952 148000 344132 148088
rect 344240 148000 344420 148088
rect 344528 148000 344708 148088
rect 344816 148000 344996 148088
rect 345104 148000 345284 148088
rect 345392 148000 345572 148088
rect 345680 148000 345860 148088
rect 346114 148000 346294 148088
rect 346402 148000 346582 148088
rect 346690 148000 346870 148088
rect 346978 148000 347158 148088
rect 347266 148000 347446 148088
rect 347554 148000 347734 148088
rect 347842 148000 348022 148088
rect 348130 148000 348310 148088
rect 348564 148000 348744 148088
rect 348852 148000 349032 148088
rect 349140 148000 349320 148088
rect 349428 148000 349608 148088
rect 349716 148000 349896 148088
rect 350004 148000 350184 148088
rect 350292 148000 350472 148088
rect 350580 148000 350760 148088
rect 351014 148000 351194 148088
rect 351302 148000 351482 148088
rect 351590 148000 351770 148088
rect 351878 148000 352058 148088
rect 352166 148000 352346 148088
rect 352454 148000 352634 148088
rect 352742 148000 352922 148088
rect 353030 148000 353210 148088
rect 353464 148000 353644 148088
rect 353752 148000 353932 148088
rect 354040 148000 354220 148088
rect 354328 148000 354508 148088
rect 354616 148000 354796 148088
rect 354904 148000 355084 148088
rect 355192 148000 355372 148088
rect 355480 148000 355660 148088
rect 355914 148000 356094 148088
rect 356202 148000 356382 148088
rect 356490 148000 356670 148088
rect 356778 148000 356958 148088
rect 357066 148000 357246 148088
rect 357354 148000 357534 148088
rect 357642 148000 357822 148088
rect 357930 148000 358110 148088
rect 358364 148000 358544 148088
rect 358652 148000 358832 148088
rect 358940 148000 359120 148088
rect 359228 148000 359408 148088
rect 359516 148000 359696 148088
rect 359804 148000 359984 148088
rect 360092 148000 360272 148088
rect 360380 148000 360560 148088
rect 360814 148000 360994 148088
rect 361102 148000 361282 148088
rect 361390 148000 361570 148088
rect 361678 148000 361858 148088
rect 361966 148000 362146 148088
rect 362254 148000 362434 148088
rect 362542 148000 362722 148088
rect 362830 148000 363010 148088
rect 363264 148000 363444 148088
rect 363552 148000 363732 148088
rect 363840 148000 364020 148088
rect 364128 148000 364308 148088
rect 364416 148000 364596 148088
rect 364704 148000 364884 148088
rect 364992 148000 365172 148088
rect 365280 148000 365460 148088
rect 365714 148000 365894 148088
rect 366002 148000 366182 148088
rect 366290 148000 366470 148088
rect 366578 148000 366758 148088
rect 366866 148000 367046 148088
rect 367154 148000 367334 148088
rect 367442 148000 367622 148088
rect 367730 148000 367910 148088
rect 243214 147784 243394 147872
rect 243502 147784 243682 147872
rect 243790 147784 243970 147872
rect 244078 147784 244258 147872
rect 244366 147784 244546 147872
rect 244654 147784 244834 147872
rect 244942 147784 245122 147872
rect 245230 147784 245410 147872
rect 245664 147784 245844 147872
rect 245952 147784 246132 147872
rect 246240 147784 246420 147872
rect 246528 147784 246708 147872
rect 246816 147784 246996 147872
rect 247104 147784 247284 147872
rect 247392 147784 247572 147872
rect 247680 147784 247860 147872
rect 248114 147784 248294 147872
rect 248402 147784 248582 147872
rect 248690 147784 248870 147872
rect 248978 147784 249158 147872
rect 249266 147784 249446 147872
rect 249554 147784 249734 147872
rect 249842 147784 250022 147872
rect 250130 147784 250310 147872
rect 250564 147784 250744 147872
rect 250852 147784 251032 147872
rect 251140 147784 251320 147872
rect 251428 147784 251608 147872
rect 251716 147784 251896 147872
rect 252004 147784 252184 147872
rect 252292 147784 252472 147872
rect 252580 147784 252760 147872
rect 253014 147784 253194 147872
rect 253302 147784 253482 147872
rect 253590 147784 253770 147872
rect 253878 147784 254058 147872
rect 254166 147784 254346 147872
rect 254454 147784 254634 147872
rect 254742 147784 254922 147872
rect 255030 147784 255210 147872
rect 255464 147784 255644 147872
rect 255752 147784 255932 147872
rect 256040 147784 256220 147872
rect 256328 147784 256508 147872
rect 256616 147784 256796 147872
rect 256904 147784 257084 147872
rect 257192 147784 257372 147872
rect 257480 147784 257660 147872
rect 257914 147784 258094 147872
rect 258202 147784 258382 147872
rect 258490 147784 258670 147872
rect 258778 147784 258958 147872
rect 259066 147784 259246 147872
rect 259354 147784 259534 147872
rect 259642 147784 259822 147872
rect 259930 147784 260110 147872
rect 260364 147784 260544 147872
rect 260652 147784 260832 147872
rect 260940 147784 261120 147872
rect 261228 147784 261408 147872
rect 261516 147784 261696 147872
rect 261804 147784 261984 147872
rect 262092 147784 262272 147872
rect 262380 147784 262560 147872
rect 262814 147784 262994 147872
rect 263102 147784 263282 147872
rect 263390 147784 263570 147872
rect 263678 147784 263858 147872
rect 263966 147784 264146 147872
rect 264254 147784 264434 147872
rect 264542 147784 264722 147872
rect 264830 147784 265010 147872
rect 265264 147784 265444 147872
rect 265552 147784 265732 147872
rect 265840 147784 266020 147872
rect 266128 147784 266308 147872
rect 266416 147784 266596 147872
rect 266704 147784 266884 147872
rect 266992 147784 267172 147872
rect 267280 147784 267460 147872
rect 267714 147784 267894 147872
rect 268002 147784 268182 147872
rect 268290 147784 268470 147872
rect 268578 147784 268758 147872
rect 268866 147784 269046 147872
rect 269154 147784 269334 147872
rect 269442 147784 269622 147872
rect 269730 147784 269910 147872
rect 270164 147784 270344 147872
rect 270452 147784 270632 147872
rect 270740 147784 270920 147872
rect 271028 147784 271208 147872
rect 271316 147784 271496 147872
rect 271604 147784 271784 147872
rect 271892 147784 272072 147872
rect 272180 147784 272360 147872
rect 272614 147784 272794 147872
rect 272902 147784 273082 147872
rect 273190 147784 273370 147872
rect 273478 147784 273658 147872
rect 273766 147784 273946 147872
rect 274054 147784 274234 147872
rect 274342 147784 274522 147872
rect 274630 147784 274810 147872
rect 275064 147784 275244 147872
rect 275352 147784 275532 147872
rect 275640 147784 275820 147872
rect 275928 147784 276108 147872
rect 276216 147784 276396 147872
rect 276504 147784 276684 147872
rect 276792 147784 276972 147872
rect 277080 147784 277260 147872
rect 277514 147784 277694 147872
rect 277802 147784 277982 147872
rect 278090 147784 278270 147872
rect 278378 147784 278558 147872
rect 278666 147784 278846 147872
rect 278954 147784 279134 147872
rect 279242 147784 279422 147872
rect 279530 147784 279710 147872
rect 279964 147784 280144 147872
rect 280252 147784 280432 147872
rect 280540 147784 280720 147872
rect 280828 147784 281008 147872
rect 281116 147784 281296 147872
rect 281404 147784 281584 147872
rect 281692 147784 281872 147872
rect 281980 147784 282160 147872
rect 282414 147784 282594 147872
rect 282702 147784 282882 147872
rect 282990 147784 283170 147872
rect 283278 147784 283458 147872
rect 283566 147784 283746 147872
rect 283854 147784 284034 147872
rect 284142 147784 284322 147872
rect 284430 147784 284610 147872
rect 284864 147784 285044 147872
rect 285152 147784 285332 147872
rect 285440 147784 285620 147872
rect 285728 147784 285908 147872
rect 286016 147784 286196 147872
rect 286304 147784 286484 147872
rect 286592 147784 286772 147872
rect 286880 147784 287060 147872
rect 287314 147784 287494 147872
rect 287602 147784 287782 147872
rect 287890 147784 288070 147872
rect 288178 147784 288358 147872
rect 288466 147784 288646 147872
rect 288754 147784 288934 147872
rect 289042 147784 289222 147872
rect 289330 147784 289510 147872
rect 289764 147784 289944 147872
rect 290052 147784 290232 147872
rect 290340 147784 290520 147872
rect 290628 147784 290808 147872
rect 290916 147784 291096 147872
rect 291204 147784 291384 147872
rect 291492 147784 291672 147872
rect 291780 147784 291960 147872
rect 292214 147784 292394 147872
rect 292502 147784 292682 147872
rect 292790 147784 292970 147872
rect 293078 147784 293258 147872
rect 293366 147784 293546 147872
rect 293654 147784 293834 147872
rect 293942 147784 294122 147872
rect 294230 147784 294410 147872
rect 294664 147784 294844 147872
rect 294952 147784 295132 147872
rect 295240 147784 295420 147872
rect 295528 147784 295708 147872
rect 295816 147784 295996 147872
rect 296104 147784 296284 147872
rect 296392 147784 296572 147872
rect 296680 147784 296860 147872
rect 297114 147784 297294 147872
rect 297402 147784 297582 147872
rect 297690 147784 297870 147872
rect 297978 147784 298158 147872
rect 298266 147784 298446 147872
rect 298554 147784 298734 147872
rect 298842 147784 299022 147872
rect 299130 147784 299310 147872
rect 299564 147784 299744 147872
rect 299852 147784 300032 147872
rect 300140 147784 300320 147872
rect 300428 147784 300608 147872
rect 300716 147784 300896 147872
rect 301004 147784 301184 147872
rect 301292 147784 301472 147872
rect 301580 147784 301760 147872
rect 302014 147784 302194 147872
rect 302302 147784 302482 147872
rect 302590 147784 302770 147872
rect 302878 147784 303058 147872
rect 303166 147784 303346 147872
rect 303454 147784 303634 147872
rect 303742 147784 303922 147872
rect 304030 147784 304210 147872
rect 304464 147784 304644 147872
rect 304752 147784 304932 147872
rect 305040 147784 305220 147872
rect 305328 147784 305508 147872
rect 305616 147784 305796 147872
rect 305904 147784 306084 147872
rect 306192 147784 306372 147872
rect 306480 147784 306660 147872
rect 306914 147784 307094 147872
rect 307202 147784 307382 147872
rect 307490 147784 307670 147872
rect 307778 147784 307958 147872
rect 308066 147784 308246 147872
rect 308354 147784 308534 147872
rect 308642 147784 308822 147872
rect 308930 147784 309110 147872
rect 309364 147784 309544 147872
rect 309652 147784 309832 147872
rect 309940 147784 310120 147872
rect 310228 147784 310408 147872
rect 310516 147784 310696 147872
rect 310804 147784 310984 147872
rect 311092 147784 311272 147872
rect 311380 147784 311560 147872
rect 311814 147784 311994 147872
rect 312102 147784 312282 147872
rect 312390 147784 312570 147872
rect 312678 147784 312858 147872
rect 312966 147784 313146 147872
rect 313254 147784 313434 147872
rect 313542 147784 313722 147872
rect 313830 147784 314010 147872
rect 314264 147784 314444 147872
rect 314552 147784 314732 147872
rect 314840 147784 315020 147872
rect 315128 147784 315308 147872
rect 315416 147784 315596 147872
rect 315704 147784 315884 147872
rect 315992 147784 316172 147872
rect 316280 147784 316460 147872
rect 316714 147784 316894 147872
rect 317002 147784 317182 147872
rect 317290 147784 317470 147872
rect 317578 147784 317758 147872
rect 317866 147784 318046 147872
rect 318154 147784 318334 147872
rect 318442 147784 318622 147872
rect 318730 147784 318910 147872
rect 319164 147784 319344 147872
rect 319452 147784 319632 147872
rect 319740 147784 319920 147872
rect 320028 147784 320208 147872
rect 320316 147784 320496 147872
rect 320604 147784 320784 147872
rect 320892 147784 321072 147872
rect 321180 147784 321360 147872
rect 321614 147784 321794 147872
rect 321902 147784 322082 147872
rect 322190 147784 322370 147872
rect 322478 147784 322658 147872
rect 322766 147784 322946 147872
rect 323054 147784 323234 147872
rect 323342 147784 323522 147872
rect 323630 147784 323810 147872
rect 324064 147784 324244 147872
rect 324352 147784 324532 147872
rect 324640 147784 324820 147872
rect 324928 147784 325108 147872
rect 325216 147784 325396 147872
rect 325504 147784 325684 147872
rect 325792 147784 325972 147872
rect 326080 147784 326260 147872
rect 326514 147784 326694 147872
rect 326802 147784 326982 147872
rect 327090 147784 327270 147872
rect 327378 147784 327558 147872
rect 327666 147784 327846 147872
rect 327954 147784 328134 147872
rect 328242 147784 328422 147872
rect 328530 147784 328710 147872
rect 328964 147784 329144 147872
rect 329252 147784 329432 147872
rect 329540 147784 329720 147872
rect 329828 147784 330008 147872
rect 330116 147784 330296 147872
rect 330404 147784 330584 147872
rect 330692 147784 330872 147872
rect 330980 147784 331160 147872
rect 331414 147784 331594 147872
rect 331702 147784 331882 147872
rect 331990 147784 332170 147872
rect 332278 147784 332458 147872
rect 332566 147784 332746 147872
rect 332854 147784 333034 147872
rect 333142 147784 333322 147872
rect 333430 147784 333610 147872
rect 333864 147784 334044 147872
rect 334152 147784 334332 147872
rect 334440 147784 334620 147872
rect 334728 147784 334908 147872
rect 335016 147784 335196 147872
rect 335304 147784 335484 147872
rect 335592 147784 335772 147872
rect 335880 147784 336060 147872
rect 336314 147784 336494 147872
rect 336602 147784 336782 147872
rect 336890 147784 337070 147872
rect 337178 147784 337358 147872
rect 337466 147784 337646 147872
rect 337754 147784 337934 147872
rect 338042 147784 338222 147872
rect 338330 147784 338510 147872
rect 338764 147784 338944 147872
rect 339052 147784 339232 147872
rect 339340 147784 339520 147872
rect 339628 147784 339808 147872
rect 339916 147784 340096 147872
rect 340204 147784 340384 147872
rect 340492 147784 340672 147872
rect 340780 147784 340960 147872
rect 341214 147784 341394 147872
rect 341502 147784 341682 147872
rect 341790 147784 341970 147872
rect 342078 147784 342258 147872
rect 342366 147784 342546 147872
rect 342654 147784 342834 147872
rect 342942 147784 343122 147872
rect 343230 147784 343410 147872
rect 343664 147784 343844 147872
rect 343952 147784 344132 147872
rect 344240 147784 344420 147872
rect 344528 147784 344708 147872
rect 344816 147784 344996 147872
rect 345104 147784 345284 147872
rect 345392 147784 345572 147872
rect 345680 147784 345860 147872
rect 346114 147784 346294 147872
rect 346402 147784 346582 147872
rect 346690 147784 346870 147872
rect 346978 147784 347158 147872
rect 347266 147784 347446 147872
rect 347554 147784 347734 147872
rect 347842 147784 348022 147872
rect 348130 147784 348310 147872
rect 348564 147784 348744 147872
rect 348852 147784 349032 147872
rect 349140 147784 349320 147872
rect 349428 147784 349608 147872
rect 349716 147784 349896 147872
rect 350004 147784 350184 147872
rect 350292 147784 350472 147872
rect 350580 147784 350760 147872
rect 351014 147784 351194 147872
rect 351302 147784 351482 147872
rect 351590 147784 351770 147872
rect 351878 147784 352058 147872
rect 352166 147784 352346 147872
rect 352454 147784 352634 147872
rect 352742 147784 352922 147872
rect 353030 147784 353210 147872
rect 353464 147784 353644 147872
rect 353752 147784 353932 147872
rect 354040 147784 354220 147872
rect 354328 147784 354508 147872
rect 354616 147784 354796 147872
rect 354904 147784 355084 147872
rect 355192 147784 355372 147872
rect 355480 147784 355660 147872
rect 355914 147784 356094 147872
rect 356202 147784 356382 147872
rect 356490 147784 356670 147872
rect 356778 147784 356958 147872
rect 357066 147784 357246 147872
rect 357354 147784 357534 147872
rect 357642 147784 357822 147872
rect 357930 147784 358110 147872
rect 358364 147784 358544 147872
rect 358652 147784 358832 147872
rect 358940 147784 359120 147872
rect 359228 147784 359408 147872
rect 359516 147784 359696 147872
rect 359804 147784 359984 147872
rect 360092 147784 360272 147872
rect 360380 147784 360560 147872
rect 360814 147784 360994 147872
rect 361102 147784 361282 147872
rect 361390 147784 361570 147872
rect 361678 147784 361858 147872
rect 361966 147784 362146 147872
rect 362254 147784 362434 147872
rect 362542 147784 362722 147872
rect 362830 147784 363010 147872
rect 363264 147784 363444 147872
rect 363552 147784 363732 147872
rect 363840 147784 364020 147872
rect 364128 147784 364308 147872
rect 364416 147784 364596 147872
rect 364704 147784 364884 147872
rect 364992 147784 365172 147872
rect 365280 147784 365460 147872
rect 365714 147784 365894 147872
rect 366002 147784 366182 147872
rect 366290 147784 366470 147872
rect 366578 147784 366758 147872
rect 366866 147784 367046 147872
rect 367154 147784 367334 147872
rect 367442 147784 367622 147872
rect 367730 147784 367910 147872
rect 243214 147308 243394 147396
rect 243502 147308 243682 147396
rect 243790 147308 243970 147396
rect 244078 147308 244258 147396
rect 244366 147308 244546 147396
rect 244654 147308 244834 147396
rect 244942 147308 245122 147396
rect 245230 147308 245410 147396
rect 245664 147308 245844 147396
rect 245952 147308 246132 147396
rect 246240 147308 246420 147396
rect 246528 147308 246708 147396
rect 246816 147308 246996 147396
rect 247104 147308 247284 147396
rect 247392 147308 247572 147396
rect 247680 147308 247860 147396
rect 248114 147308 248294 147396
rect 248402 147308 248582 147396
rect 248690 147308 248870 147396
rect 248978 147308 249158 147396
rect 249266 147308 249446 147396
rect 249554 147308 249734 147396
rect 249842 147308 250022 147396
rect 250130 147308 250310 147396
rect 250564 147308 250744 147396
rect 250852 147308 251032 147396
rect 251140 147308 251320 147396
rect 251428 147308 251608 147396
rect 251716 147308 251896 147396
rect 252004 147308 252184 147396
rect 252292 147308 252472 147396
rect 252580 147308 252760 147396
rect 253014 147308 253194 147396
rect 253302 147308 253482 147396
rect 253590 147308 253770 147396
rect 253878 147308 254058 147396
rect 254166 147308 254346 147396
rect 254454 147308 254634 147396
rect 254742 147308 254922 147396
rect 255030 147308 255210 147396
rect 255464 147308 255644 147396
rect 255752 147308 255932 147396
rect 256040 147308 256220 147396
rect 256328 147308 256508 147396
rect 256616 147308 256796 147396
rect 256904 147308 257084 147396
rect 257192 147308 257372 147396
rect 257480 147308 257660 147396
rect 257914 147308 258094 147396
rect 258202 147308 258382 147396
rect 258490 147308 258670 147396
rect 258778 147308 258958 147396
rect 259066 147308 259246 147396
rect 259354 147308 259534 147396
rect 259642 147308 259822 147396
rect 259930 147308 260110 147396
rect 260364 147308 260544 147396
rect 260652 147308 260832 147396
rect 260940 147308 261120 147396
rect 261228 147308 261408 147396
rect 261516 147308 261696 147396
rect 261804 147308 261984 147396
rect 262092 147308 262272 147396
rect 262380 147308 262560 147396
rect 262814 147308 262994 147396
rect 263102 147308 263282 147396
rect 263390 147308 263570 147396
rect 263678 147308 263858 147396
rect 263966 147308 264146 147396
rect 264254 147308 264434 147396
rect 264542 147308 264722 147396
rect 264830 147308 265010 147396
rect 265264 147308 265444 147396
rect 265552 147308 265732 147396
rect 265840 147308 266020 147396
rect 266128 147308 266308 147396
rect 266416 147308 266596 147396
rect 266704 147308 266884 147396
rect 266992 147308 267172 147396
rect 267280 147308 267460 147396
rect 267714 147308 267894 147396
rect 268002 147308 268182 147396
rect 268290 147308 268470 147396
rect 268578 147308 268758 147396
rect 268866 147308 269046 147396
rect 269154 147308 269334 147396
rect 269442 147308 269622 147396
rect 269730 147308 269910 147396
rect 270164 147308 270344 147396
rect 270452 147308 270632 147396
rect 270740 147308 270920 147396
rect 271028 147308 271208 147396
rect 271316 147308 271496 147396
rect 271604 147308 271784 147396
rect 271892 147308 272072 147396
rect 272180 147308 272360 147396
rect 272614 147308 272794 147396
rect 272902 147308 273082 147396
rect 273190 147308 273370 147396
rect 273478 147308 273658 147396
rect 273766 147308 273946 147396
rect 274054 147308 274234 147396
rect 274342 147308 274522 147396
rect 274630 147308 274810 147396
rect 275064 147308 275244 147396
rect 275352 147308 275532 147396
rect 275640 147308 275820 147396
rect 275928 147308 276108 147396
rect 276216 147308 276396 147396
rect 276504 147308 276684 147396
rect 276792 147308 276972 147396
rect 277080 147308 277260 147396
rect 277514 147308 277694 147396
rect 277802 147308 277982 147396
rect 278090 147308 278270 147396
rect 278378 147308 278558 147396
rect 278666 147308 278846 147396
rect 278954 147308 279134 147396
rect 279242 147308 279422 147396
rect 279530 147308 279710 147396
rect 279964 147308 280144 147396
rect 280252 147308 280432 147396
rect 280540 147308 280720 147396
rect 280828 147308 281008 147396
rect 281116 147308 281296 147396
rect 281404 147308 281584 147396
rect 281692 147308 281872 147396
rect 281980 147308 282160 147396
rect 282414 147308 282594 147396
rect 282702 147308 282882 147396
rect 282990 147308 283170 147396
rect 283278 147308 283458 147396
rect 283566 147308 283746 147396
rect 283854 147308 284034 147396
rect 284142 147308 284322 147396
rect 284430 147308 284610 147396
rect 284864 147308 285044 147396
rect 285152 147308 285332 147396
rect 285440 147308 285620 147396
rect 285728 147308 285908 147396
rect 286016 147308 286196 147396
rect 286304 147308 286484 147396
rect 286592 147308 286772 147396
rect 286880 147308 287060 147396
rect 287314 147308 287494 147396
rect 287602 147308 287782 147396
rect 287890 147308 288070 147396
rect 288178 147308 288358 147396
rect 288466 147308 288646 147396
rect 288754 147308 288934 147396
rect 289042 147308 289222 147396
rect 289330 147308 289510 147396
rect 289764 147308 289944 147396
rect 290052 147308 290232 147396
rect 290340 147308 290520 147396
rect 290628 147308 290808 147396
rect 290916 147308 291096 147396
rect 291204 147308 291384 147396
rect 291492 147308 291672 147396
rect 291780 147308 291960 147396
rect 292214 147308 292394 147396
rect 292502 147308 292682 147396
rect 292790 147308 292970 147396
rect 293078 147308 293258 147396
rect 293366 147308 293546 147396
rect 293654 147308 293834 147396
rect 293942 147308 294122 147396
rect 294230 147308 294410 147396
rect 294664 147308 294844 147396
rect 294952 147308 295132 147396
rect 295240 147308 295420 147396
rect 295528 147308 295708 147396
rect 295816 147308 295996 147396
rect 296104 147308 296284 147396
rect 296392 147308 296572 147396
rect 296680 147308 296860 147396
rect 297114 147308 297294 147396
rect 297402 147308 297582 147396
rect 297690 147308 297870 147396
rect 297978 147308 298158 147396
rect 298266 147308 298446 147396
rect 298554 147308 298734 147396
rect 298842 147308 299022 147396
rect 299130 147308 299310 147396
rect 299564 147308 299744 147396
rect 299852 147308 300032 147396
rect 300140 147308 300320 147396
rect 300428 147308 300608 147396
rect 300716 147308 300896 147396
rect 301004 147308 301184 147396
rect 301292 147308 301472 147396
rect 301580 147308 301760 147396
rect 302014 147308 302194 147396
rect 302302 147308 302482 147396
rect 302590 147308 302770 147396
rect 302878 147308 303058 147396
rect 303166 147308 303346 147396
rect 303454 147308 303634 147396
rect 303742 147308 303922 147396
rect 304030 147308 304210 147396
rect 304464 147308 304644 147396
rect 304752 147308 304932 147396
rect 305040 147308 305220 147396
rect 305328 147308 305508 147396
rect 305616 147308 305796 147396
rect 305904 147308 306084 147396
rect 306192 147308 306372 147396
rect 306480 147308 306660 147396
rect 306914 147308 307094 147396
rect 307202 147308 307382 147396
rect 307490 147308 307670 147396
rect 307778 147308 307958 147396
rect 308066 147308 308246 147396
rect 308354 147308 308534 147396
rect 308642 147308 308822 147396
rect 308930 147308 309110 147396
rect 309364 147308 309544 147396
rect 309652 147308 309832 147396
rect 309940 147308 310120 147396
rect 310228 147308 310408 147396
rect 310516 147308 310696 147396
rect 310804 147308 310984 147396
rect 311092 147308 311272 147396
rect 311380 147308 311560 147396
rect 311814 147308 311994 147396
rect 312102 147308 312282 147396
rect 312390 147308 312570 147396
rect 312678 147308 312858 147396
rect 312966 147308 313146 147396
rect 313254 147308 313434 147396
rect 313542 147308 313722 147396
rect 313830 147308 314010 147396
rect 314264 147308 314444 147396
rect 314552 147308 314732 147396
rect 314840 147308 315020 147396
rect 315128 147308 315308 147396
rect 315416 147308 315596 147396
rect 315704 147308 315884 147396
rect 315992 147308 316172 147396
rect 316280 147308 316460 147396
rect 316714 147308 316894 147396
rect 317002 147308 317182 147396
rect 317290 147308 317470 147396
rect 317578 147308 317758 147396
rect 317866 147308 318046 147396
rect 318154 147308 318334 147396
rect 318442 147308 318622 147396
rect 318730 147308 318910 147396
rect 319164 147308 319344 147396
rect 319452 147308 319632 147396
rect 319740 147308 319920 147396
rect 320028 147308 320208 147396
rect 320316 147308 320496 147396
rect 320604 147308 320784 147396
rect 320892 147308 321072 147396
rect 321180 147308 321360 147396
rect 321614 147308 321794 147396
rect 321902 147308 322082 147396
rect 322190 147308 322370 147396
rect 322478 147308 322658 147396
rect 322766 147308 322946 147396
rect 323054 147308 323234 147396
rect 323342 147308 323522 147396
rect 323630 147308 323810 147396
rect 324064 147308 324244 147396
rect 324352 147308 324532 147396
rect 324640 147308 324820 147396
rect 324928 147308 325108 147396
rect 325216 147308 325396 147396
rect 325504 147308 325684 147396
rect 325792 147308 325972 147396
rect 326080 147308 326260 147396
rect 326514 147308 326694 147396
rect 326802 147308 326982 147396
rect 327090 147308 327270 147396
rect 327378 147308 327558 147396
rect 327666 147308 327846 147396
rect 327954 147308 328134 147396
rect 328242 147308 328422 147396
rect 328530 147308 328710 147396
rect 328964 147308 329144 147396
rect 329252 147308 329432 147396
rect 329540 147308 329720 147396
rect 329828 147308 330008 147396
rect 330116 147308 330296 147396
rect 330404 147308 330584 147396
rect 330692 147308 330872 147396
rect 330980 147308 331160 147396
rect 331414 147308 331594 147396
rect 331702 147308 331882 147396
rect 331990 147308 332170 147396
rect 332278 147308 332458 147396
rect 332566 147308 332746 147396
rect 332854 147308 333034 147396
rect 333142 147308 333322 147396
rect 333430 147308 333610 147396
rect 333864 147308 334044 147396
rect 334152 147308 334332 147396
rect 334440 147308 334620 147396
rect 334728 147308 334908 147396
rect 335016 147308 335196 147396
rect 335304 147308 335484 147396
rect 335592 147308 335772 147396
rect 335880 147308 336060 147396
rect 336314 147308 336494 147396
rect 336602 147308 336782 147396
rect 336890 147308 337070 147396
rect 337178 147308 337358 147396
rect 337466 147308 337646 147396
rect 337754 147308 337934 147396
rect 338042 147308 338222 147396
rect 338330 147308 338510 147396
rect 338764 147308 338944 147396
rect 339052 147308 339232 147396
rect 339340 147308 339520 147396
rect 339628 147308 339808 147396
rect 339916 147308 340096 147396
rect 340204 147308 340384 147396
rect 340492 147308 340672 147396
rect 340780 147308 340960 147396
rect 341214 147308 341394 147396
rect 341502 147308 341682 147396
rect 341790 147308 341970 147396
rect 342078 147308 342258 147396
rect 342366 147308 342546 147396
rect 342654 147308 342834 147396
rect 342942 147308 343122 147396
rect 343230 147308 343410 147396
rect 343664 147308 343844 147396
rect 343952 147308 344132 147396
rect 344240 147308 344420 147396
rect 344528 147308 344708 147396
rect 344816 147308 344996 147396
rect 345104 147308 345284 147396
rect 345392 147308 345572 147396
rect 345680 147308 345860 147396
rect 346114 147308 346294 147396
rect 346402 147308 346582 147396
rect 346690 147308 346870 147396
rect 346978 147308 347158 147396
rect 347266 147308 347446 147396
rect 347554 147308 347734 147396
rect 347842 147308 348022 147396
rect 348130 147308 348310 147396
rect 348564 147308 348744 147396
rect 348852 147308 349032 147396
rect 349140 147308 349320 147396
rect 349428 147308 349608 147396
rect 349716 147308 349896 147396
rect 350004 147308 350184 147396
rect 350292 147308 350472 147396
rect 350580 147308 350760 147396
rect 351014 147308 351194 147396
rect 351302 147308 351482 147396
rect 351590 147308 351770 147396
rect 351878 147308 352058 147396
rect 352166 147308 352346 147396
rect 352454 147308 352634 147396
rect 352742 147308 352922 147396
rect 353030 147308 353210 147396
rect 353464 147308 353644 147396
rect 353752 147308 353932 147396
rect 354040 147308 354220 147396
rect 354328 147308 354508 147396
rect 354616 147308 354796 147396
rect 354904 147308 355084 147396
rect 355192 147308 355372 147396
rect 355480 147308 355660 147396
rect 355914 147308 356094 147396
rect 356202 147308 356382 147396
rect 356490 147308 356670 147396
rect 356778 147308 356958 147396
rect 357066 147308 357246 147396
rect 357354 147308 357534 147396
rect 357642 147308 357822 147396
rect 357930 147308 358110 147396
rect 358364 147308 358544 147396
rect 358652 147308 358832 147396
rect 358940 147308 359120 147396
rect 359228 147308 359408 147396
rect 359516 147308 359696 147396
rect 359804 147308 359984 147396
rect 360092 147308 360272 147396
rect 360380 147308 360560 147396
rect 360814 147308 360994 147396
rect 361102 147308 361282 147396
rect 361390 147308 361570 147396
rect 361678 147308 361858 147396
rect 361966 147308 362146 147396
rect 362254 147308 362434 147396
rect 362542 147308 362722 147396
rect 362830 147308 363010 147396
rect 363264 147308 363444 147396
rect 363552 147308 363732 147396
rect 363840 147308 364020 147396
rect 364128 147308 364308 147396
rect 364416 147308 364596 147396
rect 364704 147308 364884 147396
rect 364992 147308 365172 147396
rect 365280 147308 365460 147396
rect 365714 147308 365894 147396
rect 366002 147308 366182 147396
rect 366290 147308 366470 147396
rect 366578 147308 366758 147396
rect 366866 147308 367046 147396
rect 367154 147308 367334 147396
rect 367442 147308 367622 147396
rect 367730 147308 367910 147396
rect 243214 147092 243394 147180
rect 243502 147092 243682 147180
rect 243790 147092 243970 147180
rect 244078 147092 244258 147180
rect 244366 147092 244546 147180
rect 244654 147092 244834 147180
rect 244942 147092 245122 147180
rect 245230 147092 245410 147180
rect 245664 147092 245844 147180
rect 245952 147092 246132 147180
rect 246240 147092 246420 147180
rect 246528 147092 246708 147180
rect 246816 147092 246996 147180
rect 247104 147092 247284 147180
rect 247392 147092 247572 147180
rect 247680 147092 247860 147180
rect 248114 147092 248294 147180
rect 248402 147092 248582 147180
rect 248690 147092 248870 147180
rect 248978 147092 249158 147180
rect 249266 147092 249446 147180
rect 249554 147092 249734 147180
rect 249842 147092 250022 147180
rect 250130 147092 250310 147180
rect 250564 147092 250744 147180
rect 250852 147092 251032 147180
rect 251140 147092 251320 147180
rect 251428 147092 251608 147180
rect 251716 147092 251896 147180
rect 252004 147092 252184 147180
rect 252292 147092 252472 147180
rect 252580 147092 252760 147180
rect 253014 147092 253194 147180
rect 253302 147092 253482 147180
rect 253590 147092 253770 147180
rect 253878 147092 254058 147180
rect 254166 147092 254346 147180
rect 254454 147092 254634 147180
rect 254742 147092 254922 147180
rect 255030 147092 255210 147180
rect 255464 147092 255644 147180
rect 255752 147092 255932 147180
rect 256040 147092 256220 147180
rect 256328 147092 256508 147180
rect 256616 147092 256796 147180
rect 256904 147092 257084 147180
rect 257192 147092 257372 147180
rect 257480 147092 257660 147180
rect 257914 147092 258094 147180
rect 258202 147092 258382 147180
rect 258490 147092 258670 147180
rect 258778 147092 258958 147180
rect 259066 147092 259246 147180
rect 259354 147092 259534 147180
rect 259642 147092 259822 147180
rect 259930 147092 260110 147180
rect 260364 147092 260544 147180
rect 260652 147092 260832 147180
rect 260940 147092 261120 147180
rect 261228 147092 261408 147180
rect 261516 147092 261696 147180
rect 261804 147092 261984 147180
rect 262092 147092 262272 147180
rect 262380 147092 262560 147180
rect 262814 147092 262994 147180
rect 263102 147092 263282 147180
rect 263390 147092 263570 147180
rect 263678 147092 263858 147180
rect 263966 147092 264146 147180
rect 264254 147092 264434 147180
rect 264542 147092 264722 147180
rect 264830 147092 265010 147180
rect 265264 147092 265444 147180
rect 265552 147092 265732 147180
rect 265840 147092 266020 147180
rect 266128 147092 266308 147180
rect 266416 147092 266596 147180
rect 266704 147092 266884 147180
rect 266992 147092 267172 147180
rect 267280 147092 267460 147180
rect 267714 147092 267894 147180
rect 268002 147092 268182 147180
rect 268290 147092 268470 147180
rect 268578 147092 268758 147180
rect 268866 147092 269046 147180
rect 269154 147092 269334 147180
rect 269442 147092 269622 147180
rect 269730 147092 269910 147180
rect 270164 147092 270344 147180
rect 270452 147092 270632 147180
rect 270740 147092 270920 147180
rect 271028 147092 271208 147180
rect 271316 147092 271496 147180
rect 271604 147092 271784 147180
rect 271892 147092 272072 147180
rect 272180 147092 272360 147180
rect 272614 147092 272794 147180
rect 272902 147092 273082 147180
rect 273190 147092 273370 147180
rect 273478 147092 273658 147180
rect 273766 147092 273946 147180
rect 274054 147092 274234 147180
rect 274342 147092 274522 147180
rect 274630 147092 274810 147180
rect 275064 147092 275244 147180
rect 275352 147092 275532 147180
rect 275640 147092 275820 147180
rect 275928 147092 276108 147180
rect 276216 147092 276396 147180
rect 276504 147092 276684 147180
rect 276792 147092 276972 147180
rect 277080 147092 277260 147180
rect 277514 147092 277694 147180
rect 277802 147092 277982 147180
rect 278090 147092 278270 147180
rect 278378 147092 278558 147180
rect 278666 147092 278846 147180
rect 278954 147092 279134 147180
rect 279242 147092 279422 147180
rect 279530 147092 279710 147180
rect 279964 147092 280144 147180
rect 280252 147092 280432 147180
rect 280540 147092 280720 147180
rect 280828 147092 281008 147180
rect 281116 147092 281296 147180
rect 281404 147092 281584 147180
rect 281692 147092 281872 147180
rect 281980 147092 282160 147180
rect 282414 147092 282594 147180
rect 282702 147092 282882 147180
rect 282990 147092 283170 147180
rect 283278 147092 283458 147180
rect 283566 147092 283746 147180
rect 283854 147092 284034 147180
rect 284142 147092 284322 147180
rect 284430 147092 284610 147180
rect 284864 147092 285044 147180
rect 285152 147092 285332 147180
rect 285440 147092 285620 147180
rect 285728 147092 285908 147180
rect 286016 147092 286196 147180
rect 286304 147092 286484 147180
rect 286592 147092 286772 147180
rect 286880 147092 287060 147180
rect 287314 147092 287494 147180
rect 287602 147092 287782 147180
rect 287890 147092 288070 147180
rect 288178 147092 288358 147180
rect 288466 147092 288646 147180
rect 288754 147092 288934 147180
rect 289042 147092 289222 147180
rect 289330 147092 289510 147180
rect 289764 147092 289944 147180
rect 290052 147092 290232 147180
rect 290340 147092 290520 147180
rect 290628 147092 290808 147180
rect 290916 147092 291096 147180
rect 291204 147092 291384 147180
rect 291492 147092 291672 147180
rect 291780 147092 291960 147180
rect 292214 147092 292394 147180
rect 292502 147092 292682 147180
rect 292790 147092 292970 147180
rect 293078 147092 293258 147180
rect 293366 147092 293546 147180
rect 293654 147092 293834 147180
rect 293942 147092 294122 147180
rect 294230 147092 294410 147180
rect 294664 147092 294844 147180
rect 294952 147092 295132 147180
rect 295240 147092 295420 147180
rect 295528 147092 295708 147180
rect 295816 147092 295996 147180
rect 296104 147092 296284 147180
rect 296392 147092 296572 147180
rect 296680 147092 296860 147180
rect 297114 147092 297294 147180
rect 297402 147092 297582 147180
rect 297690 147092 297870 147180
rect 297978 147092 298158 147180
rect 298266 147092 298446 147180
rect 298554 147092 298734 147180
rect 298842 147092 299022 147180
rect 299130 147092 299310 147180
rect 299564 147092 299744 147180
rect 299852 147092 300032 147180
rect 300140 147092 300320 147180
rect 300428 147092 300608 147180
rect 300716 147092 300896 147180
rect 301004 147092 301184 147180
rect 301292 147092 301472 147180
rect 301580 147092 301760 147180
rect 302014 147092 302194 147180
rect 302302 147092 302482 147180
rect 302590 147092 302770 147180
rect 302878 147092 303058 147180
rect 303166 147092 303346 147180
rect 303454 147092 303634 147180
rect 303742 147092 303922 147180
rect 304030 147092 304210 147180
rect 304464 147092 304644 147180
rect 304752 147092 304932 147180
rect 305040 147092 305220 147180
rect 305328 147092 305508 147180
rect 305616 147092 305796 147180
rect 305904 147092 306084 147180
rect 306192 147092 306372 147180
rect 306480 147092 306660 147180
rect 306914 147092 307094 147180
rect 307202 147092 307382 147180
rect 307490 147092 307670 147180
rect 307778 147092 307958 147180
rect 308066 147092 308246 147180
rect 308354 147092 308534 147180
rect 308642 147092 308822 147180
rect 308930 147092 309110 147180
rect 309364 147092 309544 147180
rect 309652 147092 309832 147180
rect 309940 147092 310120 147180
rect 310228 147092 310408 147180
rect 310516 147092 310696 147180
rect 310804 147092 310984 147180
rect 311092 147092 311272 147180
rect 311380 147092 311560 147180
rect 311814 147092 311994 147180
rect 312102 147092 312282 147180
rect 312390 147092 312570 147180
rect 312678 147092 312858 147180
rect 312966 147092 313146 147180
rect 313254 147092 313434 147180
rect 313542 147092 313722 147180
rect 313830 147092 314010 147180
rect 314264 147092 314444 147180
rect 314552 147092 314732 147180
rect 314840 147092 315020 147180
rect 315128 147092 315308 147180
rect 315416 147092 315596 147180
rect 315704 147092 315884 147180
rect 315992 147092 316172 147180
rect 316280 147092 316460 147180
rect 316714 147092 316894 147180
rect 317002 147092 317182 147180
rect 317290 147092 317470 147180
rect 317578 147092 317758 147180
rect 317866 147092 318046 147180
rect 318154 147092 318334 147180
rect 318442 147092 318622 147180
rect 318730 147092 318910 147180
rect 319164 147092 319344 147180
rect 319452 147092 319632 147180
rect 319740 147092 319920 147180
rect 320028 147092 320208 147180
rect 320316 147092 320496 147180
rect 320604 147092 320784 147180
rect 320892 147092 321072 147180
rect 321180 147092 321360 147180
rect 321614 147092 321794 147180
rect 321902 147092 322082 147180
rect 322190 147092 322370 147180
rect 322478 147092 322658 147180
rect 322766 147092 322946 147180
rect 323054 147092 323234 147180
rect 323342 147092 323522 147180
rect 323630 147092 323810 147180
rect 324064 147092 324244 147180
rect 324352 147092 324532 147180
rect 324640 147092 324820 147180
rect 324928 147092 325108 147180
rect 325216 147092 325396 147180
rect 325504 147092 325684 147180
rect 325792 147092 325972 147180
rect 326080 147092 326260 147180
rect 326514 147092 326694 147180
rect 326802 147092 326982 147180
rect 327090 147092 327270 147180
rect 327378 147092 327558 147180
rect 327666 147092 327846 147180
rect 327954 147092 328134 147180
rect 328242 147092 328422 147180
rect 328530 147092 328710 147180
rect 328964 147092 329144 147180
rect 329252 147092 329432 147180
rect 329540 147092 329720 147180
rect 329828 147092 330008 147180
rect 330116 147092 330296 147180
rect 330404 147092 330584 147180
rect 330692 147092 330872 147180
rect 330980 147092 331160 147180
rect 331414 147092 331594 147180
rect 331702 147092 331882 147180
rect 331990 147092 332170 147180
rect 332278 147092 332458 147180
rect 332566 147092 332746 147180
rect 332854 147092 333034 147180
rect 333142 147092 333322 147180
rect 333430 147092 333610 147180
rect 333864 147092 334044 147180
rect 334152 147092 334332 147180
rect 334440 147092 334620 147180
rect 334728 147092 334908 147180
rect 335016 147092 335196 147180
rect 335304 147092 335484 147180
rect 335592 147092 335772 147180
rect 335880 147092 336060 147180
rect 336314 147092 336494 147180
rect 336602 147092 336782 147180
rect 336890 147092 337070 147180
rect 337178 147092 337358 147180
rect 337466 147092 337646 147180
rect 337754 147092 337934 147180
rect 338042 147092 338222 147180
rect 338330 147092 338510 147180
rect 338764 147092 338944 147180
rect 339052 147092 339232 147180
rect 339340 147092 339520 147180
rect 339628 147092 339808 147180
rect 339916 147092 340096 147180
rect 340204 147092 340384 147180
rect 340492 147092 340672 147180
rect 340780 147092 340960 147180
rect 341214 147092 341394 147180
rect 341502 147092 341682 147180
rect 341790 147092 341970 147180
rect 342078 147092 342258 147180
rect 342366 147092 342546 147180
rect 342654 147092 342834 147180
rect 342942 147092 343122 147180
rect 343230 147092 343410 147180
rect 343664 147092 343844 147180
rect 343952 147092 344132 147180
rect 344240 147092 344420 147180
rect 344528 147092 344708 147180
rect 344816 147092 344996 147180
rect 345104 147092 345284 147180
rect 345392 147092 345572 147180
rect 345680 147092 345860 147180
rect 346114 147092 346294 147180
rect 346402 147092 346582 147180
rect 346690 147092 346870 147180
rect 346978 147092 347158 147180
rect 347266 147092 347446 147180
rect 347554 147092 347734 147180
rect 347842 147092 348022 147180
rect 348130 147092 348310 147180
rect 348564 147092 348744 147180
rect 348852 147092 349032 147180
rect 349140 147092 349320 147180
rect 349428 147092 349608 147180
rect 349716 147092 349896 147180
rect 350004 147092 350184 147180
rect 350292 147092 350472 147180
rect 350580 147092 350760 147180
rect 351014 147092 351194 147180
rect 351302 147092 351482 147180
rect 351590 147092 351770 147180
rect 351878 147092 352058 147180
rect 352166 147092 352346 147180
rect 352454 147092 352634 147180
rect 352742 147092 352922 147180
rect 353030 147092 353210 147180
rect 353464 147092 353644 147180
rect 353752 147092 353932 147180
rect 354040 147092 354220 147180
rect 354328 147092 354508 147180
rect 354616 147092 354796 147180
rect 354904 147092 355084 147180
rect 355192 147092 355372 147180
rect 355480 147092 355660 147180
rect 355914 147092 356094 147180
rect 356202 147092 356382 147180
rect 356490 147092 356670 147180
rect 356778 147092 356958 147180
rect 357066 147092 357246 147180
rect 357354 147092 357534 147180
rect 357642 147092 357822 147180
rect 357930 147092 358110 147180
rect 358364 147092 358544 147180
rect 358652 147092 358832 147180
rect 358940 147092 359120 147180
rect 359228 147092 359408 147180
rect 359516 147092 359696 147180
rect 359804 147092 359984 147180
rect 360092 147092 360272 147180
rect 360380 147092 360560 147180
rect 360814 147092 360994 147180
rect 361102 147092 361282 147180
rect 361390 147092 361570 147180
rect 361678 147092 361858 147180
rect 361966 147092 362146 147180
rect 362254 147092 362434 147180
rect 362542 147092 362722 147180
rect 362830 147092 363010 147180
rect 363264 147092 363444 147180
rect 363552 147092 363732 147180
rect 363840 147092 364020 147180
rect 364128 147092 364308 147180
rect 364416 147092 364596 147180
rect 364704 147092 364884 147180
rect 364992 147092 365172 147180
rect 365280 147092 365460 147180
rect 365714 147092 365894 147180
rect 366002 147092 366182 147180
rect 366290 147092 366470 147180
rect 366578 147092 366758 147180
rect 366866 147092 367046 147180
rect 367154 147092 367334 147180
rect 367442 147092 367622 147180
rect 367730 147092 367910 147180
rect 243214 146616 243394 146704
rect 243502 146616 243682 146704
rect 243790 146616 243970 146704
rect 244078 146616 244258 146704
rect 244366 146616 244546 146704
rect 244654 146616 244834 146704
rect 244942 146616 245122 146704
rect 245230 146616 245410 146704
rect 245664 146616 245844 146704
rect 245952 146616 246132 146704
rect 246240 146616 246420 146704
rect 246528 146616 246708 146704
rect 246816 146616 246996 146704
rect 247104 146616 247284 146704
rect 247392 146616 247572 146704
rect 247680 146616 247860 146704
rect 248114 146616 248294 146704
rect 248402 146616 248582 146704
rect 248690 146616 248870 146704
rect 248978 146616 249158 146704
rect 249266 146616 249446 146704
rect 249554 146616 249734 146704
rect 249842 146616 250022 146704
rect 250130 146616 250310 146704
rect 250564 146616 250744 146704
rect 250852 146616 251032 146704
rect 251140 146616 251320 146704
rect 251428 146616 251608 146704
rect 251716 146616 251896 146704
rect 252004 146616 252184 146704
rect 252292 146616 252472 146704
rect 252580 146616 252760 146704
rect 253014 146616 253194 146704
rect 253302 146616 253482 146704
rect 253590 146616 253770 146704
rect 253878 146616 254058 146704
rect 254166 146616 254346 146704
rect 254454 146616 254634 146704
rect 254742 146616 254922 146704
rect 255030 146616 255210 146704
rect 255464 146616 255644 146704
rect 255752 146616 255932 146704
rect 256040 146616 256220 146704
rect 256328 146616 256508 146704
rect 256616 146616 256796 146704
rect 256904 146616 257084 146704
rect 257192 146616 257372 146704
rect 257480 146616 257660 146704
rect 257914 146616 258094 146704
rect 258202 146616 258382 146704
rect 258490 146616 258670 146704
rect 258778 146616 258958 146704
rect 259066 146616 259246 146704
rect 259354 146616 259534 146704
rect 259642 146616 259822 146704
rect 259930 146616 260110 146704
rect 260364 146616 260544 146704
rect 260652 146616 260832 146704
rect 260940 146616 261120 146704
rect 261228 146616 261408 146704
rect 261516 146616 261696 146704
rect 261804 146616 261984 146704
rect 262092 146616 262272 146704
rect 262380 146616 262560 146704
rect 262814 146616 262994 146704
rect 263102 146616 263282 146704
rect 263390 146616 263570 146704
rect 263678 146616 263858 146704
rect 263966 146616 264146 146704
rect 264254 146616 264434 146704
rect 264542 146616 264722 146704
rect 264830 146616 265010 146704
rect 265264 146616 265444 146704
rect 265552 146616 265732 146704
rect 265840 146616 266020 146704
rect 266128 146616 266308 146704
rect 266416 146616 266596 146704
rect 266704 146616 266884 146704
rect 266992 146616 267172 146704
rect 267280 146616 267460 146704
rect 267714 146616 267894 146704
rect 268002 146616 268182 146704
rect 268290 146616 268470 146704
rect 268578 146616 268758 146704
rect 268866 146616 269046 146704
rect 269154 146616 269334 146704
rect 269442 146616 269622 146704
rect 269730 146616 269910 146704
rect 270164 146616 270344 146704
rect 270452 146616 270632 146704
rect 270740 146616 270920 146704
rect 271028 146616 271208 146704
rect 271316 146616 271496 146704
rect 271604 146616 271784 146704
rect 271892 146616 272072 146704
rect 272180 146616 272360 146704
rect 272614 146616 272794 146704
rect 272902 146616 273082 146704
rect 273190 146616 273370 146704
rect 273478 146616 273658 146704
rect 273766 146616 273946 146704
rect 274054 146616 274234 146704
rect 274342 146616 274522 146704
rect 274630 146616 274810 146704
rect 275064 146616 275244 146704
rect 275352 146616 275532 146704
rect 275640 146616 275820 146704
rect 275928 146616 276108 146704
rect 276216 146616 276396 146704
rect 276504 146616 276684 146704
rect 276792 146616 276972 146704
rect 277080 146616 277260 146704
rect 277514 146616 277694 146704
rect 277802 146616 277982 146704
rect 278090 146616 278270 146704
rect 278378 146616 278558 146704
rect 278666 146616 278846 146704
rect 278954 146616 279134 146704
rect 279242 146616 279422 146704
rect 279530 146616 279710 146704
rect 279964 146616 280144 146704
rect 280252 146616 280432 146704
rect 280540 146616 280720 146704
rect 280828 146616 281008 146704
rect 281116 146616 281296 146704
rect 281404 146616 281584 146704
rect 281692 146616 281872 146704
rect 281980 146616 282160 146704
rect 282414 146616 282594 146704
rect 282702 146616 282882 146704
rect 282990 146616 283170 146704
rect 283278 146616 283458 146704
rect 283566 146616 283746 146704
rect 283854 146616 284034 146704
rect 284142 146616 284322 146704
rect 284430 146616 284610 146704
rect 284864 146616 285044 146704
rect 285152 146616 285332 146704
rect 285440 146616 285620 146704
rect 285728 146616 285908 146704
rect 286016 146616 286196 146704
rect 286304 146616 286484 146704
rect 286592 146616 286772 146704
rect 286880 146616 287060 146704
rect 287314 146616 287494 146704
rect 287602 146616 287782 146704
rect 287890 146616 288070 146704
rect 288178 146616 288358 146704
rect 288466 146616 288646 146704
rect 288754 146616 288934 146704
rect 289042 146616 289222 146704
rect 289330 146616 289510 146704
rect 289764 146616 289944 146704
rect 290052 146616 290232 146704
rect 290340 146616 290520 146704
rect 290628 146616 290808 146704
rect 290916 146616 291096 146704
rect 291204 146616 291384 146704
rect 291492 146616 291672 146704
rect 291780 146616 291960 146704
rect 292214 146616 292394 146704
rect 292502 146616 292682 146704
rect 292790 146616 292970 146704
rect 293078 146616 293258 146704
rect 293366 146616 293546 146704
rect 293654 146616 293834 146704
rect 293942 146616 294122 146704
rect 294230 146616 294410 146704
rect 294664 146616 294844 146704
rect 294952 146616 295132 146704
rect 295240 146616 295420 146704
rect 295528 146616 295708 146704
rect 295816 146616 295996 146704
rect 296104 146616 296284 146704
rect 296392 146616 296572 146704
rect 296680 146616 296860 146704
rect 297114 146616 297294 146704
rect 297402 146616 297582 146704
rect 297690 146616 297870 146704
rect 297978 146616 298158 146704
rect 298266 146616 298446 146704
rect 298554 146616 298734 146704
rect 298842 146616 299022 146704
rect 299130 146616 299310 146704
rect 299564 146616 299744 146704
rect 299852 146616 300032 146704
rect 300140 146616 300320 146704
rect 300428 146616 300608 146704
rect 300716 146616 300896 146704
rect 301004 146616 301184 146704
rect 301292 146616 301472 146704
rect 301580 146616 301760 146704
rect 302014 146616 302194 146704
rect 302302 146616 302482 146704
rect 302590 146616 302770 146704
rect 302878 146616 303058 146704
rect 303166 146616 303346 146704
rect 303454 146616 303634 146704
rect 303742 146616 303922 146704
rect 304030 146616 304210 146704
rect 304464 146616 304644 146704
rect 304752 146616 304932 146704
rect 305040 146616 305220 146704
rect 305328 146616 305508 146704
rect 305616 146616 305796 146704
rect 305904 146616 306084 146704
rect 306192 146616 306372 146704
rect 306480 146616 306660 146704
rect 306914 146616 307094 146704
rect 307202 146616 307382 146704
rect 307490 146616 307670 146704
rect 307778 146616 307958 146704
rect 308066 146616 308246 146704
rect 308354 146616 308534 146704
rect 308642 146616 308822 146704
rect 308930 146616 309110 146704
rect 309364 146616 309544 146704
rect 309652 146616 309832 146704
rect 309940 146616 310120 146704
rect 310228 146616 310408 146704
rect 310516 146616 310696 146704
rect 310804 146616 310984 146704
rect 311092 146616 311272 146704
rect 311380 146616 311560 146704
rect 311814 146616 311994 146704
rect 312102 146616 312282 146704
rect 312390 146616 312570 146704
rect 312678 146616 312858 146704
rect 312966 146616 313146 146704
rect 313254 146616 313434 146704
rect 313542 146616 313722 146704
rect 313830 146616 314010 146704
rect 314264 146616 314444 146704
rect 314552 146616 314732 146704
rect 314840 146616 315020 146704
rect 315128 146616 315308 146704
rect 315416 146616 315596 146704
rect 315704 146616 315884 146704
rect 315992 146616 316172 146704
rect 316280 146616 316460 146704
rect 316714 146616 316894 146704
rect 317002 146616 317182 146704
rect 317290 146616 317470 146704
rect 317578 146616 317758 146704
rect 317866 146616 318046 146704
rect 318154 146616 318334 146704
rect 318442 146616 318622 146704
rect 318730 146616 318910 146704
rect 319164 146616 319344 146704
rect 319452 146616 319632 146704
rect 319740 146616 319920 146704
rect 320028 146616 320208 146704
rect 320316 146616 320496 146704
rect 320604 146616 320784 146704
rect 320892 146616 321072 146704
rect 321180 146616 321360 146704
rect 321614 146616 321794 146704
rect 321902 146616 322082 146704
rect 322190 146616 322370 146704
rect 322478 146616 322658 146704
rect 322766 146616 322946 146704
rect 323054 146616 323234 146704
rect 323342 146616 323522 146704
rect 323630 146616 323810 146704
rect 324064 146616 324244 146704
rect 324352 146616 324532 146704
rect 324640 146616 324820 146704
rect 324928 146616 325108 146704
rect 325216 146616 325396 146704
rect 325504 146616 325684 146704
rect 325792 146616 325972 146704
rect 326080 146616 326260 146704
rect 326514 146616 326694 146704
rect 326802 146616 326982 146704
rect 327090 146616 327270 146704
rect 327378 146616 327558 146704
rect 327666 146616 327846 146704
rect 327954 146616 328134 146704
rect 328242 146616 328422 146704
rect 328530 146616 328710 146704
rect 328964 146616 329144 146704
rect 329252 146616 329432 146704
rect 329540 146616 329720 146704
rect 329828 146616 330008 146704
rect 330116 146616 330296 146704
rect 330404 146616 330584 146704
rect 330692 146616 330872 146704
rect 330980 146616 331160 146704
rect 331414 146616 331594 146704
rect 331702 146616 331882 146704
rect 331990 146616 332170 146704
rect 332278 146616 332458 146704
rect 332566 146616 332746 146704
rect 332854 146616 333034 146704
rect 333142 146616 333322 146704
rect 333430 146616 333610 146704
rect 333864 146616 334044 146704
rect 334152 146616 334332 146704
rect 334440 146616 334620 146704
rect 334728 146616 334908 146704
rect 335016 146616 335196 146704
rect 335304 146616 335484 146704
rect 335592 146616 335772 146704
rect 335880 146616 336060 146704
rect 336314 146616 336494 146704
rect 336602 146616 336782 146704
rect 336890 146616 337070 146704
rect 337178 146616 337358 146704
rect 337466 146616 337646 146704
rect 337754 146616 337934 146704
rect 338042 146616 338222 146704
rect 338330 146616 338510 146704
rect 338764 146616 338944 146704
rect 339052 146616 339232 146704
rect 339340 146616 339520 146704
rect 339628 146616 339808 146704
rect 339916 146616 340096 146704
rect 340204 146616 340384 146704
rect 340492 146616 340672 146704
rect 340780 146616 340960 146704
rect 341214 146616 341394 146704
rect 341502 146616 341682 146704
rect 341790 146616 341970 146704
rect 342078 146616 342258 146704
rect 342366 146616 342546 146704
rect 342654 146616 342834 146704
rect 342942 146616 343122 146704
rect 343230 146616 343410 146704
rect 343664 146616 343844 146704
rect 343952 146616 344132 146704
rect 344240 146616 344420 146704
rect 344528 146616 344708 146704
rect 344816 146616 344996 146704
rect 345104 146616 345284 146704
rect 345392 146616 345572 146704
rect 345680 146616 345860 146704
rect 346114 146616 346294 146704
rect 346402 146616 346582 146704
rect 346690 146616 346870 146704
rect 346978 146616 347158 146704
rect 347266 146616 347446 146704
rect 347554 146616 347734 146704
rect 347842 146616 348022 146704
rect 348130 146616 348310 146704
rect 348564 146616 348744 146704
rect 348852 146616 349032 146704
rect 349140 146616 349320 146704
rect 349428 146616 349608 146704
rect 349716 146616 349896 146704
rect 350004 146616 350184 146704
rect 350292 146616 350472 146704
rect 350580 146616 350760 146704
rect 351014 146616 351194 146704
rect 351302 146616 351482 146704
rect 351590 146616 351770 146704
rect 351878 146616 352058 146704
rect 352166 146616 352346 146704
rect 352454 146616 352634 146704
rect 352742 146616 352922 146704
rect 353030 146616 353210 146704
rect 353464 146616 353644 146704
rect 353752 146616 353932 146704
rect 354040 146616 354220 146704
rect 354328 146616 354508 146704
rect 354616 146616 354796 146704
rect 354904 146616 355084 146704
rect 355192 146616 355372 146704
rect 355480 146616 355660 146704
rect 355914 146616 356094 146704
rect 356202 146616 356382 146704
rect 356490 146616 356670 146704
rect 356778 146616 356958 146704
rect 357066 146616 357246 146704
rect 357354 146616 357534 146704
rect 357642 146616 357822 146704
rect 357930 146616 358110 146704
rect 358364 146616 358544 146704
rect 358652 146616 358832 146704
rect 358940 146616 359120 146704
rect 359228 146616 359408 146704
rect 359516 146616 359696 146704
rect 359804 146616 359984 146704
rect 360092 146616 360272 146704
rect 360380 146616 360560 146704
rect 360814 146616 360994 146704
rect 361102 146616 361282 146704
rect 361390 146616 361570 146704
rect 361678 146616 361858 146704
rect 361966 146616 362146 146704
rect 362254 146616 362434 146704
rect 362542 146616 362722 146704
rect 362830 146616 363010 146704
rect 363264 146616 363444 146704
rect 363552 146616 363732 146704
rect 363840 146616 364020 146704
rect 364128 146616 364308 146704
rect 364416 146616 364596 146704
rect 364704 146616 364884 146704
rect 364992 146616 365172 146704
rect 365280 146616 365460 146704
rect 365714 146616 365894 146704
rect 366002 146616 366182 146704
rect 366290 146616 366470 146704
rect 366578 146616 366758 146704
rect 366866 146616 367046 146704
rect 367154 146616 367334 146704
rect 367442 146616 367622 146704
rect 367730 146616 367910 146704
rect 243214 146400 243394 146488
rect 243502 146400 243682 146488
rect 243790 146400 243970 146488
rect 244078 146400 244258 146488
rect 244366 146400 244546 146488
rect 244654 146400 244834 146488
rect 244942 146400 245122 146488
rect 245230 146400 245410 146488
rect 245664 146400 245844 146488
rect 245952 146400 246132 146488
rect 246240 146400 246420 146488
rect 246528 146400 246708 146488
rect 246816 146400 246996 146488
rect 247104 146400 247284 146488
rect 247392 146400 247572 146488
rect 247680 146400 247860 146488
rect 248114 146400 248294 146488
rect 248402 146400 248582 146488
rect 248690 146400 248870 146488
rect 248978 146400 249158 146488
rect 249266 146400 249446 146488
rect 249554 146400 249734 146488
rect 249842 146400 250022 146488
rect 250130 146400 250310 146488
rect 250564 146400 250744 146488
rect 250852 146400 251032 146488
rect 251140 146400 251320 146488
rect 251428 146400 251608 146488
rect 251716 146400 251896 146488
rect 252004 146400 252184 146488
rect 252292 146400 252472 146488
rect 252580 146400 252760 146488
rect 253014 146400 253194 146488
rect 253302 146400 253482 146488
rect 253590 146400 253770 146488
rect 253878 146400 254058 146488
rect 254166 146400 254346 146488
rect 254454 146400 254634 146488
rect 254742 146400 254922 146488
rect 255030 146400 255210 146488
rect 255464 146400 255644 146488
rect 255752 146400 255932 146488
rect 256040 146400 256220 146488
rect 256328 146400 256508 146488
rect 256616 146400 256796 146488
rect 256904 146400 257084 146488
rect 257192 146400 257372 146488
rect 257480 146400 257660 146488
rect 257914 146400 258094 146488
rect 258202 146400 258382 146488
rect 258490 146400 258670 146488
rect 258778 146400 258958 146488
rect 259066 146400 259246 146488
rect 259354 146400 259534 146488
rect 259642 146400 259822 146488
rect 259930 146400 260110 146488
rect 260364 146400 260544 146488
rect 260652 146400 260832 146488
rect 260940 146400 261120 146488
rect 261228 146400 261408 146488
rect 261516 146400 261696 146488
rect 261804 146400 261984 146488
rect 262092 146400 262272 146488
rect 262380 146400 262560 146488
rect 262814 146400 262994 146488
rect 263102 146400 263282 146488
rect 263390 146400 263570 146488
rect 263678 146400 263858 146488
rect 263966 146400 264146 146488
rect 264254 146400 264434 146488
rect 264542 146400 264722 146488
rect 264830 146400 265010 146488
rect 265264 146400 265444 146488
rect 265552 146400 265732 146488
rect 265840 146400 266020 146488
rect 266128 146400 266308 146488
rect 266416 146400 266596 146488
rect 266704 146400 266884 146488
rect 266992 146400 267172 146488
rect 267280 146400 267460 146488
rect 267714 146400 267894 146488
rect 268002 146400 268182 146488
rect 268290 146400 268470 146488
rect 268578 146400 268758 146488
rect 268866 146400 269046 146488
rect 269154 146400 269334 146488
rect 269442 146400 269622 146488
rect 269730 146400 269910 146488
rect 270164 146400 270344 146488
rect 270452 146400 270632 146488
rect 270740 146400 270920 146488
rect 271028 146400 271208 146488
rect 271316 146400 271496 146488
rect 271604 146400 271784 146488
rect 271892 146400 272072 146488
rect 272180 146400 272360 146488
rect 272614 146400 272794 146488
rect 272902 146400 273082 146488
rect 273190 146400 273370 146488
rect 273478 146400 273658 146488
rect 273766 146400 273946 146488
rect 274054 146400 274234 146488
rect 274342 146400 274522 146488
rect 274630 146400 274810 146488
rect 275064 146400 275244 146488
rect 275352 146400 275532 146488
rect 275640 146400 275820 146488
rect 275928 146400 276108 146488
rect 276216 146400 276396 146488
rect 276504 146400 276684 146488
rect 276792 146400 276972 146488
rect 277080 146400 277260 146488
rect 277514 146400 277694 146488
rect 277802 146400 277982 146488
rect 278090 146400 278270 146488
rect 278378 146400 278558 146488
rect 278666 146400 278846 146488
rect 278954 146400 279134 146488
rect 279242 146400 279422 146488
rect 279530 146400 279710 146488
rect 279964 146400 280144 146488
rect 280252 146400 280432 146488
rect 280540 146400 280720 146488
rect 280828 146400 281008 146488
rect 281116 146400 281296 146488
rect 281404 146400 281584 146488
rect 281692 146400 281872 146488
rect 281980 146400 282160 146488
rect 282414 146400 282594 146488
rect 282702 146400 282882 146488
rect 282990 146400 283170 146488
rect 283278 146400 283458 146488
rect 283566 146400 283746 146488
rect 283854 146400 284034 146488
rect 284142 146400 284322 146488
rect 284430 146400 284610 146488
rect 284864 146400 285044 146488
rect 285152 146400 285332 146488
rect 285440 146400 285620 146488
rect 285728 146400 285908 146488
rect 286016 146400 286196 146488
rect 286304 146400 286484 146488
rect 286592 146400 286772 146488
rect 286880 146400 287060 146488
rect 287314 146400 287494 146488
rect 287602 146400 287782 146488
rect 287890 146400 288070 146488
rect 288178 146400 288358 146488
rect 288466 146400 288646 146488
rect 288754 146400 288934 146488
rect 289042 146400 289222 146488
rect 289330 146400 289510 146488
rect 289764 146400 289944 146488
rect 290052 146400 290232 146488
rect 290340 146400 290520 146488
rect 290628 146400 290808 146488
rect 290916 146400 291096 146488
rect 291204 146400 291384 146488
rect 291492 146400 291672 146488
rect 291780 146400 291960 146488
rect 292214 146400 292394 146488
rect 292502 146400 292682 146488
rect 292790 146400 292970 146488
rect 293078 146400 293258 146488
rect 293366 146400 293546 146488
rect 293654 146400 293834 146488
rect 293942 146400 294122 146488
rect 294230 146400 294410 146488
rect 294664 146400 294844 146488
rect 294952 146400 295132 146488
rect 295240 146400 295420 146488
rect 295528 146400 295708 146488
rect 295816 146400 295996 146488
rect 296104 146400 296284 146488
rect 296392 146400 296572 146488
rect 296680 146400 296860 146488
rect 297114 146400 297294 146488
rect 297402 146400 297582 146488
rect 297690 146400 297870 146488
rect 297978 146400 298158 146488
rect 298266 146400 298446 146488
rect 298554 146400 298734 146488
rect 298842 146400 299022 146488
rect 299130 146400 299310 146488
rect 299564 146400 299744 146488
rect 299852 146400 300032 146488
rect 300140 146400 300320 146488
rect 300428 146400 300608 146488
rect 300716 146400 300896 146488
rect 301004 146400 301184 146488
rect 301292 146400 301472 146488
rect 301580 146400 301760 146488
rect 302014 146400 302194 146488
rect 302302 146400 302482 146488
rect 302590 146400 302770 146488
rect 302878 146400 303058 146488
rect 303166 146400 303346 146488
rect 303454 146400 303634 146488
rect 303742 146400 303922 146488
rect 304030 146400 304210 146488
rect 304464 146400 304644 146488
rect 304752 146400 304932 146488
rect 305040 146400 305220 146488
rect 305328 146400 305508 146488
rect 305616 146400 305796 146488
rect 305904 146400 306084 146488
rect 306192 146400 306372 146488
rect 306480 146400 306660 146488
rect 306914 146400 307094 146488
rect 307202 146400 307382 146488
rect 307490 146400 307670 146488
rect 307778 146400 307958 146488
rect 308066 146400 308246 146488
rect 308354 146400 308534 146488
rect 308642 146400 308822 146488
rect 308930 146400 309110 146488
rect 309364 146400 309544 146488
rect 309652 146400 309832 146488
rect 309940 146400 310120 146488
rect 310228 146400 310408 146488
rect 310516 146400 310696 146488
rect 310804 146400 310984 146488
rect 311092 146400 311272 146488
rect 311380 146400 311560 146488
rect 311814 146400 311994 146488
rect 312102 146400 312282 146488
rect 312390 146400 312570 146488
rect 312678 146400 312858 146488
rect 312966 146400 313146 146488
rect 313254 146400 313434 146488
rect 313542 146400 313722 146488
rect 313830 146400 314010 146488
rect 314264 146400 314444 146488
rect 314552 146400 314732 146488
rect 314840 146400 315020 146488
rect 315128 146400 315308 146488
rect 315416 146400 315596 146488
rect 315704 146400 315884 146488
rect 315992 146400 316172 146488
rect 316280 146400 316460 146488
rect 316714 146400 316894 146488
rect 317002 146400 317182 146488
rect 317290 146400 317470 146488
rect 317578 146400 317758 146488
rect 317866 146400 318046 146488
rect 318154 146400 318334 146488
rect 318442 146400 318622 146488
rect 318730 146400 318910 146488
rect 319164 146400 319344 146488
rect 319452 146400 319632 146488
rect 319740 146400 319920 146488
rect 320028 146400 320208 146488
rect 320316 146400 320496 146488
rect 320604 146400 320784 146488
rect 320892 146400 321072 146488
rect 321180 146400 321360 146488
rect 321614 146400 321794 146488
rect 321902 146400 322082 146488
rect 322190 146400 322370 146488
rect 322478 146400 322658 146488
rect 322766 146400 322946 146488
rect 323054 146400 323234 146488
rect 323342 146400 323522 146488
rect 323630 146400 323810 146488
rect 324064 146400 324244 146488
rect 324352 146400 324532 146488
rect 324640 146400 324820 146488
rect 324928 146400 325108 146488
rect 325216 146400 325396 146488
rect 325504 146400 325684 146488
rect 325792 146400 325972 146488
rect 326080 146400 326260 146488
rect 326514 146400 326694 146488
rect 326802 146400 326982 146488
rect 327090 146400 327270 146488
rect 327378 146400 327558 146488
rect 327666 146400 327846 146488
rect 327954 146400 328134 146488
rect 328242 146400 328422 146488
rect 328530 146400 328710 146488
rect 328964 146400 329144 146488
rect 329252 146400 329432 146488
rect 329540 146400 329720 146488
rect 329828 146400 330008 146488
rect 330116 146400 330296 146488
rect 330404 146400 330584 146488
rect 330692 146400 330872 146488
rect 330980 146400 331160 146488
rect 331414 146400 331594 146488
rect 331702 146400 331882 146488
rect 331990 146400 332170 146488
rect 332278 146400 332458 146488
rect 332566 146400 332746 146488
rect 332854 146400 333034 146488
rect 333142 146400 333322 146488
rect 333430 146400 333610 146488
rect 333864 146400 334044 146488
rect 334152 146400 334332 146488
rect 334440 146400 334620 146488
rect 334728 146400 334908 146488
rect 335016 146400 335196 146488
rect 335304 146400 335484 146488
rect 335592 146400 335772 146488
rect 335880 146400 336060 146488
rect 336314 146400 336494 146488
rect 336602 146400 336782 146488
rect 336890 146400 337070 146488
rect 337178 146400 337358 146488
rect 337466 146400 337646 146488
rect 337754 146400 337934 146488
rect 338042 146400 338222 146488
rect 338330 146400 338510 146488
rect 338764 146400 338944 146488
rect 339052 146400 339232 146488
rect 339340 146400 339520 146488
rect 339628 146400 339808 146488
rect 339916 146400 340096 146488
rect 340204 146400 340384 146488
rect 340492 146400 340672 146488
rect 340780 146400 340960 146488
rect 341214 146400 341394 146488
rect 341502 146400 341682 146488
rect 341790 146400 341970 146488
rect 342078 146400 342258 146488
rect 342366 146400 342546 146488
rect 342654 146400 342834 146488
rect 342942 146400 343122 146488
rect 343230 146400 343410 146488
rect 343664 146400 343844 146488
rect 343952 146400 344132 146488
rect 344240 146400 344420 146488
rect 344528 146400 344708 146488
rect 344816 146400 344996 146488
rect 345104 146400 345284 146488
rect 345392 146400 345572 146488
rect 345680 146400 345860 146488
rect 346114 146400 346294 146488
rect 346402 146400 346582 146488
rect 346690 146400 346870 146488
rect 346978 146400 347158 146488
rect 347266 146400 347446 146488
rect 347554 146400 347734 146488
rect 347842 146400 348022 146488
rect 348130 146400 348310 146488
rect 348564 146400 348744 146488
rect 348852 146400 349032 146488
rect 349140 146400 349320 146488
rect 349428 146400 349608 146488
rect 349716 146400 349896 146488
rect 350004 146400 350184 146488
rect 350292 146400 350472 146488
rect 350580 146400 350760 146488
rect 351014 146400 351194 146488
rect 351302 146400 351482 146488
rect 351590 146400 351770 146488
rect 351878 146400 352058 146488
rect 352166 146400 352346 146488
rect 352454 146400 352634 146488
rect 352742 146400 352922 146488
rect 353030 146400 353210 146488
rect 353464 146400 353644 146488
rect 353752 146400 353932 146488
rect 354040 146400 354220 146488
rect 354328 146400 354508 146488
rect 354616 146400 354796 146488
rect 354904 146400 355084 146488
rect 355192 146400 355372 146488
rect 355480 146400 355660 146488
rect 355914 146400 356094 146488
rect 356202 146400 356382 146488
rect 356490 146400 356670 146488
rect 356778 146400 356958 146488
rect 357066 146400 357246 146488
rect 357354 146400 357534 146488
rect 357642 146400 357822 146488
rect 357930 146400 358110 146488
rect 358364 146400 358544 146488
rect 358652 146400 358832 146488
rect 358940 146400 359120 146488
rect 359228 146400 359408 146488
rect 359516 146400 359696 146488
rect 359804 146400 359984 146488
rect 360092 146400 360272 146488
rect 360380 146400 360560 146488
rect 360814 146400 360994 146488
rect 361102 146400 361282 146488
rect 361390 146400 361570 146488
rect 361678 146400 361858 146488
rect 361966 146400 362146 146488
rect 362254 146400 362434 146488
rect 362542 146400 362722 146488
rect 362830 146400 363010 146488
rect 363264 146400 363444 146488
rect 363552 146400 363732 146488
rect 363840 146400 364020 146488
rect 364128 146400 364308 146488
rect 364416 146400 364596 146488
rect 364704 146400 364884 146488
rect 364992 146400 365172 146488
rect 365280 146400 365460 146488
rect 365714 146400 365894 146488
rect 366002 146400 366182 146488
rect 366290 146400 366470 146488
rect 366578 146400 366758 146488
rect 366866 146400 367046 146488
rect 367154 146400 367334 146488
rect 367442 146400 367622 146488
rect 367730 146400 367910 146488
rect 243214 145924 243394 146012
rect 243502 145924 243682 146012
rect 243790 145924 243970 146012
rect 244078 145924 244258 146012
rect 244366 145924 244546 146012
rect 244654 145924 244834 146012
rect 244942 145924 245122 146012
rect 245230 145924 245410 146012
rect 245664 145924 245844 146012
rect 245952 145924 246132 146012
rect 246240 145924 246420 146012
rect 246528 145924 246708 146012
rect 246816 145924 246996 146012
rect 247104 145924 247284 146012
rect 247392 145924 247572 146012
rect 247680 145924 247860 146012
rect 248114 145924 248294 146012
rect 248402 145924 248582 146012
rect 248690 145924 248870 146012
rect 248978 145924 249158 146012
rect 249266 145924 249446 146012
rect 249554 145924 249734 146012
rect 249842 145924 250022 146012
rect 250130 145924 250310 146012
rect 250564 145924 250744 146012
rect 250852 145924 251032 146012
rect 251140 145924 251320 146012
rect 251428 145924 251608 146012
rect 251716 145924 251896 146012
rect 252004 145924 252184 146012
rect 252292 145924 252472 146012
rect 252580 145924 252760 146012
rect 253014 145924 253194 146012
rect 253302 145924 253482 146012
rect 253590 145924 253770 146012
rect 253878 145924 254058 146012
rect 254166 145924 254346 146012
rect 254454 145924 254634 146012
rect 254742 145924 254922 146012
rect 255030 145924 255210 146012
rect 255464 145924 255644 146012
rect 255752 145924 255932 146012
rect 256040 145924 256220 146012
rect 256328 145924 256508 146012
rect 256616 145924 256796 146012
rect 256904 145924 257084 146012
rect 257192 145924 257372 146012
rect 257480 145924 257660 146012
rect 257914 145924 258094 146012
rect 258202 145924 258382 146012
rect 258490 145924 258670 146012
rect 258778 145924 258958 146012
rect 259066 145924 259246 146012
rect 259354 145924 259534 146012
rect 259642 145924 259822 146012
rect 259930 145924 260110 146012
rect 260364 145924 260544 146012
rect 260652 145924 260832 146012
rect 260940 145924 261120 146012
rect 261228 145924 261408 146012
rect 261516 145924 261696 146012
rect 261804 145924 261984 146012
rect 262092 145924 262272 146012
rect 262380 145924 262560 146012
rect 262814 145924 262994 146012
rect 263102 145924 263282 146012
rect 263390 145924 263570 146012
rect 263678 145924 263858 146012
rect 263966 145924 264146 146012
rect 264254 145924 264434 146012
rect 264542 145924 264722 146012
rect 264830 145924 265010 146012
rect 265264 145924 265444 146012
rect 265552 145924 265732 146012
rect 265840 145924 266020 146012
rect 266128 145924 266308 146012
rect 266416 145924 266596 146012
rect 266704 145924 266884 146012
rect 266992 145924 267172 146012
rect 267280 145924 267460 146012
rect 267714 145924 267894 146012
rect 268002 145924 268182 146012
rect 268290 145924 268470 146012
rect 268578 145924 268758 146012
rect 268866 145924 269046 146012
rect 269154 145924 269334 146012
rect 269442 145924 269622 146012
rect 269730 145924 269910 146012
rect 270164 145924 270344 146012
rect 270452 145924 270632 146012
rect 270740 145924 270920 146012
rect 271028 145924 271208 146012
rect 271316 145924 271496 146012
rect 271604 145924 271784 146012
rect 271892 145924 272072 146012
rect 272180 145924 272360 146012
rect 272614 145924 272794 146012
rect 272902 145924 273082 146012
rect 273190 145924 273370 146012
rect 273478 145924 273658 146012
rect 273766 145924 273946 146012
rect 274054 145924 274234 146012
rect 274342 145924 274522 146012
rect 274630 145924 274810 146012
rect 275064 145924 275244 146012
rect 275352 145924 275532 146012
rect 275640 145924 275820 146012
rect 275928 145924 276108 146012
rect 276216 145924 276396 146012
rect 276504 145924 276684 146012
rect 276792 145924 276972 146012
rect 277080 145924 277260 146012
rect 277514 145924 277694 146012
rect 277802 145924 277982 146012
rect 278090 145924 278270 146012
rect 278378 145924 278558 146012
rect 278666 145924 278846 146012
rect 278954 145924 279134 146012
rect 279242 145924 279422 146012
rect 279530 145924 279710 146012
rect 279964 145924 280144 146012
rect 280252 145924 280432 146012
rect 280540 145924 280720 146012
rect 280828 145924 281008 146012
rect 281116 145924 281296 146012
rect 281404 145924 281584 146012
rect 281692 145924 281872 146012
rect 281980 145924 282160 146012
rect 282414 145924 282594 146012
rect 282702 145924 282882 146012
rect 282990 145924 283170 146012
rect 283278 145924 283458 146012
rect 283566 145924 283746 146012
rect 283854 145924 284034 146012
rect 284142 145924 284322 146012
rect 284430 145924 284610 146012
rect 284864 145924 285044 146012
rect 285152 145924 285332 146012
rect 285440 145924 285620 146012
rect 285728 145924 285908 146012
rect 286016 145924 286196 146012
rect 286304 145924 286484 146012
rect 286592 145924 286772 146012
rect 286880 145924 287060 146012
rect 287314 145924 287494 146012
rect 287602 145924 287782 146012
rect 287890 145924 288070 146012
rect 288178 145924 288358 146012
rect 288466 145924 288646 146012
rect 288754 145924 288934 146012
rect 289042 145924 289222 146012
rect 289330 145924 289510 146012
rect 289764 145924 289944 146012
rect 290052 145924 290232 146012
rect 290340 145924 290520 146012
rect 290628 145924 290808 146012
rect 290916 145924 291096 146012
rect 291204 145924 291384 146012
rect 291492 145924 291672 146012
rect 291780 145924 291960 146012
rect 292214 145924 292394 146012
rect 292502 145924 292682 146012
rect 292790 145924 292970 146012
rect 293078 145924 293258 146012
rect 293366 145924 293546 146012
rect 293654 145924 293834 146012
rect 293942 145924 294122 146012
rect 294230 145924 294410 146012
rect 294664 145924 294844 146012
rect 294952 145924 295132 146012
rect 295240 145924 295420 146012
rect 295528 145924 295708 146012
rect 295816 145924 295996 146012
rect 296104 145924 296284 146012
rect 296392 145924 296572 146012
rect 296680 145924 296860 146012
rect 297114 145924 297294 146012
rect 297402 145924 297582 146012
rect 297690 145924 297870 146012
rect 297978 145924 298158 146012
rect 298266 145924 298446 146012
rect 298554 145924 298734 146012
rect 298842 145924 299022 146012
rect 299130 145924 299310 146012
rect 299564 145924 299744 146012
rect 299852 145924 300032 146012
rect 300140 145924 300320 146012
rect 300428 145924 300608 146012
rect 300716 145924 300896 146012
rect 301004 145924 301184 146012
rect 301292 145924 301472 146012
rect 301580 145924 301760 146012
rect 302014 145924 302194 146012
rect 302302 145924 302482 146012
rect 302590 145924 302770 146012
rect 302878 145924 303058 146012
rect 303166 145924 303346 146012
rect 303454 145924 303634 146012
rect 303742 145924 303922 146012
rect 304030 145924 304210 146012
rect 304464 145924 304644 146012
rect 304752 145924 304932 146012
rect 305040 145924 305220 146012
rect 305328 145924 305508 146012
rect 305616 145924 305796 146012
rect 305904 145924 306084 146012
rect 306192 145924 306372 146012
rect 306480 145924 306660 146012
rect 306914 145924 307094 146012
rect 307202 145924 307382 146012
rect 307490 145924 307670 146012
rect 307778 145924 307958 146012
rect 308066 145924 308246 146012
rect 308354 145924 308534 146012
rect 308642 145924 308822 146012
rect 308930 145924 309110 146012
rect 309364 145924 309544 146012
rect 309652 145924 309832 146012
rect 309940 145924 310120 146012
rect 310228 145924 310408 146012
rect 310516 145924 310696 146012
rect 310804 145924 310984 146012
rect 311092 145924 311272 146012
rect 311380 145924 311560 146012
rect 311814 145924 311994 146012
rect 312102 145924 312282 146012
rect 312390 145924 312570 146012
rect 312678 145924 312858 146012
rect 312966 145924 313146 146012
rect 313254 145924 313434 146012
rect 313542 145924 313722 146012
rect 313830 145924 314010 146012
rect 314264 145924 314444 146012
rect 314552 145924 314732 146012
rect 314840 145924 315020 146012
rect 315128 145924 315308 146012
rect 315416 145924 315596 146012
rect 315704 145924 315884 146012
rect 315992 145924 316172 146012
rect 316280 145924 316460 146012
rect 316714 145924 316894 146012
rect 317002 145924 317182 146012
rect 317290 145924 317470 146012
rect 317578 145924 317758 146012
rect 317866 145924 318046 146012
rect 318154 145924 318334 146012
rect 318442 145924 318622 146012
rect 318730 145924 318910 146012
rect 319164 145924 319344 146012
rect 319452 145924 319632 146012
rect 319740 145924 319920 146012
rect 320028 145924 320208 146012
rect 320316 145924 320496 146012
rect 320604 145924 320784 146012
rect 320892 145924 321072 146012
rect 321180 145924 321360 146012
rect 321614 145924 321794 146012
rect 321902 145924 322082 146012
rect 322190 145924 322370 146012
rect 322478 145924 322658 146012
rect 322766 145924 322946 146012
rect 323054 145924 323234 146012
rect 323342 145924 323522 146012
rect 323630 145924 323810 146012
rect 324064 145924 324244 146012
rect 324352 145924 324532 146012
rect 324640 145924 324820 146012
rect 324928 145924 325108 146012
rect 325216 145924 325396 146012
rect 325504 145924 325684 146012
rect 325792 145924 325972 146012
rect 326080 145924 326260 146012
rect 326514 145924 326694 146012
rect 326802 145924 326982 146012
rect 327090 145924 327270 146012
rect 327378 145924 327558 146012
rect 327666 145924 327846 146012
rect 327954 145924 328134 146012
rect 328242 145924 328422 146012
rect 328530 145924 328710 146012
rect 328964 145924 329144 146012
rect 329252 145924 329432 146012
rect 329540 145924 329720 146012
rect 329828 145924 330008 146012
rect 330116 145924 330296 146012
rect 330404 145924 330584 146012
rect 330692 145924 330872 146012
rect 330980 145924 331160 146012
rect 331414 145924 331594 146012
rect 331702 145924 331882 146012
rect 331990 145924 332170 146012
rect 332278 145924 332458 146012
rect 332566 145924 332746 146012
rect 332854 145924 333034 146012
rect 333142 145924 333322 146012
rect 333430 145924 333610 146012
rect 333864 145924 334044 146012
rect 334152 145924 334332 146012
rect 334440 145924 334620 146012
rect 334728 145924 334908 146012
rect 335016 145924 335196 146012
rect 335304 145924 335484 146012
rect 335592 145924 335772 146012
rect 335880 145924 336060 146012
rect 336314 145924 336494 146012
rect 336602 145924 336782 146012
rect 336890 145924 337070 146012
rect 337178 145924 337358 146012
rect 337466 145924 337646 146012
rect 337754 145924 337934 146012
rect 338042 145924 338222 146012
rect 338330 145924 338510 146012
rect 338764 145924 338944 146012
rect 339052 145924 339232 146012
rect 339340 145924 339520 146012
rect 339628 145924 339808 146012
rect 339916 145924 340096 146012
rect 340204 145924 340384 146012
rect 340492 145924 340672 146012
rect 340780 145924 340960 146012
rect 341214 145924 341394 146012
rect 341502 145924 341682 146012
rect 341790 145924 341970 146012
rect 342078 145924 342258 146012
rect 342366 145924 342546 146012
rect 342654 145924 342834 146012
rect 342942 145924 343122 146012
rect 343230 145924 343410 146012
rect 343664 145924 343844 146012
rect 343952 145924 344132 146012
rect 344240 145924 344420 146012
rect 344528 145924 344708 146012
rect 344816 145924 344996 146012
rect 345104 145924 345284 146012
rect 345392 145924 345572 146012
rect 345680 145924 345860 146012
rect 346114 145924 346294 146012
rect 346402 145924 346582 146012
rect 346690 145924 346870 146012
rect 346978 145924 347158 146012
rect 347266 145924 347446 146012
rect 347554 145924 347734 146012
rect 347842 145924 348022 146012
rect 348130 145924 348310 146012
rect 348564 145924 348744 146012
rect 348852 145924 349032 146012
rect 349140 145924 349320 146012
rect 349428 145924 349608 146012
rect 349716 145924 349896 146012
rect 350004 145924 350184 146012
rect 350292 145924 350472 146012
rect 350580 145924 350760 146012
rect 351014 145924 351194 146012
rect 351302 145924 351482 146012
rect 351590 145924 351770 146012
rect 351878 145924 352058 146012
rect 352166 145924 352346 146012
rect 352454 145924 352634 146012
rect 352742 145924 352922 146012
rect 353030 145924 353210 146012
rect 353464 145924 353644 146012
rect 353752 145924 353932 146012
rect 354040 145924 354220 146012
rect 354328 145924 354508 146012
rect 354616 145924 354796 146012
rect 354904 145924 355084 146012
rect 355192 145924 355372 146012
rect 355480 145924 355660 146012
rect 355914 145924 356094 146012
rect 356202 145924 356382 146012
rect 356490 145924 356670 146012
rect 356778 145924 356958 146012
rect 357066 145924 357246 146012
rect 357354 145924 357534 146012
rect 357642 145924 357822 146012
rect 357930 145924 358110 146012
rect 358364 145924 358544 146012
rect 358652 145924 358832 146012
rect 358940 145924 359120 146012
rect 359228 145924 359408 146012
rect 359516 145924 359696 146012
rect 359804 145924 359984 146012
rect 360092 145924 360272 146012
rect 360380 145924 360560 146012
rect 360814 145924 360994 146012
rect 361102 145924 361282 146012
rect 361390 145924 361570 146012
rect 361678 145924 361858 146012
rect 361966 145924 362146 146012
rect 362254 145924 362434 146012
rect 362542 145924 362722 146012
rect 362830 145924 363010 146012
rect 363264 145924 363444 146012
rect 363552 145924 363732 146012
rect 363840 145924 364020 146012
rect 364128 145924 364308 146012
rect 364416 145924 364596 146012
rect 364704 145924 364884 146012
rect 364992 145924 365172 146012
rect 365280 145924 365460 146012
rect 365714 145924 365894 146012
rect 366002 145924 366182 146012
rect 366290 145924 366470 146012
rect 366578 145924 366758 146012
rect 366866 145924 367046 146012
rect 367154 145924 367334 146012
rect 367442 145924 367622 146012
rect 367730 145924 367910 146012
rect 243214 145450 243394 145538
rect 243502 145450 243682 145538
rect 243790 145450 243970 145538
rect 244078 145450 244258 145538
rect 244366 145450 244546 145538
rect 244654 145450 244834 145538
rect 244942 145450 245122 145538
rect 245230 145450 245410 145538
rect 245664 145450 245844 145538
rect 245952 145450 246132 145538
rect 246240 145450 246420 145538
rect 246528 145450 246708 145538
rect 246816 145450 246996 145538
rect 247104 145450 247284 145538
rect 247392 145450 247572 145538
rect 247680 145450 247860 145538
rect 248114 145450 248294 145538
rect 248402 145450 248582 145538
rect 248690 145450 248870 145538
rect 248978 145450 249158 145538
rect 249266 145450 249446 145538
rect 249554 145450 249734 145538
rect 249842 145450 250022 145538
rect 250130 145450 250310 145538
rect 250564 145450 250744 145538
rect 250852 145450 251032 145538
rect 251140 145450 251320 145538
rect 251428 145450 251608 145538
rect 251716 145450 251896 145538
rect 252004 145450 252184 145538
rect 252292 145450 252472 145538
rect 252580 145450 252760 145538
rect 253014 145450 253194 145538
rect 253302 145450 253482 145538
rect 253590 145450 253770 145538
rect 253878 145450 254058 145538
rect 254166 145450 254346 145538
rect 254454 145450 254634 145538
rect 254742 145450 254922 145538
rect 255030 145450 255210 145538
rect 255464 145450 255644 145538
rect 255752 145450 255932 145538
rect 256040 145450 256220 145538
rect 256328 145450 256508 145538
rect 256616 145450 256796 145538
rect 256904 145450 257084 145538
rect 257192 145450 257372 145538
rect 257480 145450 257660 145538
rect 257914 145450 258094 145538
rect 258202 145450 258382 145538
rect 258490 145450 258670 145538
rect 258778 145450 258958 145538
rect 259066 145450 259246 145538
rect 259354 145450 259534 145538
rect 259642 145450 259822 145538
rect 259930 145450 260110 145538
rect 260364 145450 260544 145538
rect 260652 145450 260832 145538
rect 260940 145450 261120 145538
rect 261228 145450 261408 145538
rect 261516 145450 261696 145538
rect 261804 145450 261984 145538
rect 262092 145450 262272 145538
rect 262380 145450 262560 145538
rect 262814 145450 262994 145538
rect 263102 145450 263282 145538
rect 263390 145450 263570 145538
rect 263678 145450 263858 145538
rect 263966 145450 264146 145538
rect 264254 145450 264434 145538
rect 264542 145450 264722 145538
rect 264830 145450 265010 145538
rect 265264 145450 265444 145538
rect 265552 145450 265732 145538
rect 265840 145450 266020 145538
rect 266128 145450 266308 145538
rect 266416 145450 266596 145538
rect 266704 145450 266884 145538
rect 266992 145450 267172 145538
rect 267280 145450 267460 145538
rect 267714 145450 267894 145538
rect 268002 145450 268182 145538
rect 268290 145450 268470 145538
rect 268578 145450 268758 145538
rect 268866 145450 269046 145538
rect 269154 145450 269334 145538
rect 269442 145450 269622 145538
rect 269730 145450 269910 145538
rect 270164 145450 270344 145538
rect 270452 145450 270632 145538
rect 270740 145450 270920 145538
rect 271028 145450 271208 145538
rect 271316 145450 271496 145538
rect 271604 145450 271784 145538
rect 271892 145450 272072 145538
rect 272180 145450 272360 145538
rect 272614 145450 272794 145538
rect 272902 145450 273082 145538
rect 273190 145450 273370 145538
rect 273478 145450 273658 145538
rect 273766 145450 273946 145538
rect 274054 145450 274234 145538
rect 274342 145450 274522 145538
rect 274630 145450 274810 145538
rect 275064 145450 275244 145538
rect 275352 145450 275532 145538
rect 275640 145450 275820 145538
rect 275928 145450 276108 145538
rect 276216 145450 276396 145538
rect 276504 145450 276684 145538
rect 276792 145450 276972 145538
rect 277080 145450 277260 145538
rect 277514 145450 277694 145538
rect 277802 145450 277982 145538
rect 278090 145450 278270 145538
rect 278378 145450 278558 145538
rect 278666 145450 278846 145538
rect 278954 145450 279134 145538
rect 279242 145450 279422 145538
rect 279530 145450 279710 145538
rect 279964 145450 280144 145538
rect 280252 145450 280432 145538
rect 280540 145450 280720 145538
rect 280828 145450 281008 145538
rect 281116 145450 281296 145538
rect 281404 145450 281584 145538
rect 281692 145450 281872 145538
rect 281980 145450 282160 145538
rect 282414 145450 282594 145538
rect 282702 145450 282882 145538
rect 282990 145450 283170 145538
rect 283278 145450 283458 145538
rect 283566 145450 283746 145538
rect 283854 145450 284034 145538
rect 284142 145450 284322 145538
rect 284430 145450 284610 145538
rect 284864 145450 285044 145538
rect 285152 145450 285332 145538
rect 285440 145450 285620 145538
rect 285728 145450 285908 145538
rect 286016 145450 286196 145538
rect 286304 145450 286484 145538
rect 286592 145450 286772 145538
rect 286880 145450 287060 145538
rect 287314 145450 287494 145538
rect 287602 145450 287782 145538
rect 287890 145450 288070 145538
rect 288178 145450 288358 145538
rect 288466 145450 288646 145538
rect 288754 145450 288934 145538
rect 289042 145450 289222 145538
rect 289330 145450 289510 145538
rect 289764 145450 289944 145538
rect 290052 145450 290232 145538
rect 290340 145450 290520 145538
rect 290628 145450 290808 145538
rect 290916 145450 291096 145538
rect 291204 145450 291384 145538
rect 291492 145450 291672 145538
rect 291780 145450 291960 145538
rect 292214 145450 292394 145538
rect 292502 145450 292682 145538
rect 292790 145450 292970 145538
rect 293078 145450 293258 145538
rect 293366 145450 293546 145538
rect 293654 145450 293834 145538
rect 293942 145450 294122 145538
rect 294230 145450 294410 145538
rect 294664 145450 294844 145538
rect 294952 145450 295132 145538
rect 295240 145450 295420 145538
rect 295528 145450 295708 145538
rect 295816 145450 295996 145538
rect 296104 145450 296284 145538
rect 296392 145450 296572 145538
rect 296680 145450 296860 145538
rect 297114 145450 297294 145538
rect 297402 145450 297582 145538
rect 297690 145450 297870 145538
rect 297978 145450 298158 145538
rect 298266 145450 298446 145538
rect 298554 145450 298734 145538
rect 298842 145450 299022 145538
rect 299130 145450 299310 145538
rect 299564 145450 299744 145538
rect 299852 145450 300032 145538
rect 300140 145450 300320 145538
rect 300428 145450 300608 145538
rect 300716 145450 300896 145538
rect 301004 145450 301184 145538
rect 301292 145450 301472 145538
rect 301580 145450 301760 145538
rect 302014 145450 302194 145538
rect 302302 145450 302482 145538
rect 302590 145450 302770 145538
rect 302878 145450 303058 145538
rect 303166 145450 303346 145538
rect 303454 145450 303634 145538
rect 303742 145450 303922 145538
rect 304030 145450 304210 145538
rect 304464 145450 304644 145538
rect 304752 145450 304932 145538
rect 305040 145450 305220 145538
rect 305328 145450 305508 145538
rect 305616 145450 305796 145538
rect 305904 145450 306084 145538
rect 306192 145450 306372 145538
rect 306480 145450 306660 145538
rect 306914 145450 307094 145538
rect 307202 145450 307382 145538
rect 307490 145450 307670 145538
rect 307778 145450 307958 145538
rect 308066 145450 308246 145538
rect 308354 145450 308534 145538
rect 308642 145450 308822 145538
rect 308930 145450 309110 145538
rect 309364 145450 309544 145538
rect 309652 145450 309832 145538
rect 309940 145450 310120 145538
rect 310228 145450 310408 145538
rect 310516 145450 310696 145538
rect 310804 145450 310984 145538
rect 311092 145450 311272 145538
rect 311380 145450 311560 145538
rect 311814 145450 311994 145538
rect 312102 145450 312282 145538
rect 312390 145450 312570 145538
rect 312678 145450 312858 145538
rect 312966 145450 313146 145538
rect 313254 145450 313434 145538
rect 313542 145450 313722 145538
rect 313830 145450 314010 145538
rect 314264 145450 314444 145538
rect 314552 145450 314732 145538
rect 314840 145450 315020 145538
rect 315128 145450 315308 145538
rect 315416 145450 315596 145538
rect 315704 145450 315884 145538
rect 315992 145450 316172 145538
rect 316280 145450 316460 145538
rect 316714 145450 316894 145538
rect 317002 145450 317182 145538
rect 317290 145450 317470 145538
rect 317578 145450 317758 145538
rect 317866 145450 318046 145538
rect 318154 145450 318334 145538
rect 318442 145450 318622 145538
rect 318730 145450 318910 145538
rect 319164 145450 319344 145538
rect 319452 145450 319632 145538
rect 319740 145450 319920 145538
rect 320028 145450 320208 145538
rect 320316 145450 320496 145538
rect 320604 145450 320784 145538
rect 320892 145450 321072 145538
rect 321180 145450 321360 145538
rect 321614 145450 321794 145538
rect 321902 145450 322082 145538
rect 322190 145450 322370 145538
rect 322478 145450 322658 145538
rect 322766 145450 322946 145538
rect 323054 145450 323234 145538
rect 323342 145450 323522 145538
rect 323630 145450 323810 145538
rect 324064 145450 324244 145538
rect 324352 145450 324532 145538
rect 324640 145450 324820 145538
rect 324928 145450 325108 145538
rect 325216 145450 325396 145538
rect 325504 145450 325684 145538
rect 325792 145450 325972 145538
rect 326080 145450 326260 145538
rect 326514 145450 326694 145538
rect 326802 145450 326982 145538
rect 327090 145450 327270 145538
rect 327378 145450 327558 145538
rect 327666 145450 327846 145538
rect 327954 145450 328134 145538
rect 328242 145450 328422 145538
rect 328530 145450 328710 145538
rect 328964 145450 329144 145538
rect 329252 145450 329432 145538
rect 329540 145450 329720 145538
rect 329828 145450 330008 145538
rect 330116 145450 330296 145538
rect 330404 145450 330584 145538
rect 330692 145450 330872 145538
rect 330980 145450 331160 145538
rect 331414 145450 331594 145538
rect 331702 145450 331882 145538
rect 331990 145450 332170 145538
rect 332278 145450 332458 145538
rect 332566 145450 332746 145538
rect 332854 145450 333034 145538
rect 333142 145450 333322 145538
rect 333430 145450 333610 145538
rect 333864 145450 334044 145538
rect 334152 145450 334332 145538
rect 334440 145450 334620 145538
rect 334728 145450 334908 145538
rect 335016 145450 335196 145538
rect 335304 145450 335484 145538
rect 335592 145450 335772 145538
rect 335880 145450 336060 145538
rect 336314 145450 336494 145538
rect 336602 145450 336782 145538
rect 336890 145450 337070 145538
rect 337178 145450 337358 145538
rect 337466 145450 337646 145538
rect 337754 145450 337934 145538
rect 338042 145450 338222 145538
rect 338330 145450 338510 145538
rect 338764 145450 338944 145538
rect 339052 145450 339232 145538
rect 339340 145450 339520 145538
rect 339628 145450 339808 145538
rect 339916 145450 340096 145538
rect 340204 145450 340384 145538
rect 340492 145450 340672 145538
rect 340780 145450 340960 145538
rect 341214 145450 341394 145538
rect 341502 145450 341682 145538
rect 341790 145450 341970 145538
rect 342078 145450 342258 145538
rect 342366 145450 342546 145538
rect 342654 145450 342834 145538
rect 342942 145450 343122 145538
rect 343230 145450 343410 145538
rect 343664 145450 343844 145538
rect 343952 145450 344132 145538
rect 344240 145450 344420 145538
rect 344528 145450 344708 145538
rect 344816 145450 344996 145538
rect 345104 145450 345284 145538
rect 345392 145450 345572 145538
rect 345680 145450 345860 145538
rect 346114 145450 346294 145538
rect 346402 145450 346582 145538
rect 346690 145450 346870 145538
rect 346978 145450 347158 145538
rect 347266 145450 347446 145538
rect 347554 145450 347734 145538
rect 347842 145450 348022 145538
rect 348130 145450 348310 145538
rect 348564 145450 348744 145538
rect 348852 145450 349032 145538
rect 349140 145450 349320 145538
rect 349428 145450 349608 145538
rect 349716 145450 349896 145538
rect 350004 145450 350184 145538
rect 350292 145450 350472 145538
rect 350580 145450 350760 145538
rect 351014 145450 351194 145538
rect 351302 145450 351482 145538
rect 351590 145450 351770 145538
rect 351878 145450 352058 145538
rect 352166 145450 352346 145538
rect 352454 145450 352634 145538
rect 352742 145450 352922 145538
rect 353030 145450 353210 145538
rect 353464 145450 353644 145538
rect 353752 145450 353932 145538
rect 354040 145450 354220 145538
rect 354328 145450 354508 145538
rect 354616 145450 354796 145538
rect 354904 145450 355084 145538
rect 355192 145450 355372 145538
rect 355480 145450 355660 145538
rect 355914 145450 356094 145538
rect 356202 145450 356382 145538
rect 356490 145450 356670 145538
rect 356778 145450 356958 145538
rect 357066 145450 357246 145538
rect 357354 145450 357534 145538
rect 357642 145450 357822 145538
rect 357930 145450 358110 145538
rect 358364 145450 358544 145538
rect 358652 145450 358832 145538
rect 358940 145450 359120 145538
rect 359228 145450 359408 145538
rect 359516 145450 359696 145538
rect 359804 145450 359984 145538
rect 360092 145450 360272 145538
rect 360380 145450 360560 145538
rect 360814 145450 360994 145538
rect 361102 145450 361282 145538
rect 361390 145450 361570 145538
rect 361678 145450 361858 145538
rect 361966 145450 362146 145538
rect 362254 145450 362434 145538
rect 362542 145450 362722 145538
rect 362830 145450 363010 145538
rect 363264 145450 363444 145538
rect 363552 145450 363732 145538
rect 363840 145450 364020 145538
rect 364128 145450 364308 145538
rect 364416 145450 364596 145538
rect 364704 145450 364884 145538
rect 364992 145450 365172 145538
rect 365280 145450 365460 145538
rect 365714 145450 365894 145538
rect 366002 145450 366182 145538
rect 366290 145450 366470 145538
rect 366578 145450 366758 145538
rect 366866 145450 367046 145538
rect 367154 145450 367334 145538
rect 367442 145450 367622 145538
rect 367730 145450 367910 145538
rect 243214 144974 243394 145062
rect 243502 144974 243682 145062
rect 243790 144974 243970 145062
rect 244078 144974 244258 145062
rect 244366 144974 244546 145062
rect 244654 144974 244834 145062
rect 244942 144974 245122 145062
rect 245230 144974 245410 145062
rect 245664 144974 245844 145062
rect 245952 144974 246132 145062
rect 246240 144974 246420 145062
rect 246528 144974 246708 145062
rect 246816 144974 246996 145062
rect 247104 144974 247284 145062
rect 247392 144974 247572 145062
rect 247680 144974 247860 145062
rect 248114 144974 248294 145062
rect 248402 144974 248582 145062
rect 248690 144974 248870 145062
rect 248978 144974 249158 145062
rect 249266 144974 249446 145062
rect 249554 144974 249734 145062
rect 249842 144974 250022 145062
rect 250130 144974 250310 145062
rect 250564 144974 250744 145062
rect 250852 144974 251032 145062
rect 251140 144974 251320 145062
rect 251428 144974 251608 145062
rect 251716 144974 251896 145062
rect 252004 144974 252184 145062
rect 252292 144974 252472 145062
rect 252580 144974 252760 145062
rect 253014 144974 253194 145062
rect 253302 144974 253482 145062
rect 253590 144974 253770 145062
rect 253878 144974 254058 145062
rect 254166 144974 254346 145062
rect 254454 144974 254634 145062
rect 254742 144974 254922 145062
rect 255030 144974 255210 145062
rect 255464 144974 255644 145062
rect 255752 144974 255932 145062
rect 256040 144974 256220 145062
rect 256328 144974 256508 145062
rect 256616 144974 256796 145062
rect 256904 144974 257084 145062
rect 257192 144974 257372 145062
rect 257480 144974 257660 145062
rect 257914 144974 258094 145062
rect 258202 144974 258382 145062
rect 258490 144974 258670 145062
rect 258778 144974 258958 145062
rect 259066 144974 259246 145062
rect 259354 144974 259534 145062
rect 259642 144974 259822 145062
rect 259930 144974 260110 145062
rect 260364 144974 260544 145062
rect 260652 144974 260832 145062
rect 260940 144974 261120 145062
rect 261228 144974 261408 145062
rect 261516 144974 261696 145062
rect 261804 144974 261984 145062
rect 262092 144974 262272 145062
rect 262380 144974 262560 145062
rect 262814 144974 262994 145062
rect 263102 144974 263282 145062
rect 263390 144974 263570 145062
rect 263678 144974 263858 145062
rect 263966 144974 264146 145062
rect 264254 144974 264434 145062
rect 264542 144974 264722 145062
rect 264830 144974 265010 145062
rect 265264 144974 265444 145062
rect 265552 144974 265732 145062
rect 265840 144974 266020 145062
rect 266128 144974 266308 145062
rect 266416 144974 266596 145062
rect 266704 144974 266884 145062
rect 266992 144974 267172 145062
rect 267280 144974 267460 145062
rect 267714 144974 267894 145062
rect 268002 144974 268182 145062
rect 268290 144974 268470 145062
rect 268578 144974 268758 145062
rect 268866 144974 269046 145062
rect 269154 144974 269334 145062
rect 269442 144974 269622 145062
rect 269730 144974 269910 145062
rect 270164 144974 270344 145062
rect 270452 144974 270632 145062
rect 270740 144974 270920 145062
rect 271028 144974 271208 145062
rect 271316 144974 271496 145062
rect 271604 144974 271784 145062
rect 271892 144974 272072 145062
rect 272180 144974 272360 145062
rect 272614 144974 272794 145062
rect 272902 144974 273082 145062
rect 273190 144974 273370 145062
rect 273478 144974 273658 145062
rect 273766 144974 273946 145062
rect 274054 144974 274234 145062
rect 274342 144974 274522 145062
rect 274630 144974 274810 145062
rect 275064 144974 275244 145062
rect 275352 144974 275532 145062
rect 275640 144974 275820 145062
rect 275928 144974 276108 145062
rect 276216 144974 276396 145062
rect 276504 144974 276684 145062
rect 276792 144974 276972 145062
rect 277080 144974 277260 145062
rect 277514 144974 277694 145062
rect 277802 144974 277982 145062
rect 278090 144974 278270 145062
rect 278378 144974 278558 145062
rect 278666 144974 278846 145062
rect 278954 144974 279134 145062
rect 279242 144974 279422 145062
rect 279530 144974 279710 145062
rect 279964 144974 280144 145062
rect 280252 144974 280432 145062
rect 280540 144974 280720 145062
rect 280828 144974 281008 145062
rect 281116 144974 281296 145062
rect 281404 144974 281584 145062
rect 281692 144974 281872 145062
rect 281980 144974 282160 145062
rect 282414 144974 282594 145062
rect 282702 144974 282882 145062
rect 282990 144974 283170 145062
rect 283278 144974 283458 145062
rect 283566 144974 283746 145062
rect 283854 144974 284034 145062
rect 284142 144974 284322 145062
rect 284430 144974 284610 145062
rect 284864 144974 285044 145062
rect 285152 144974 285332 145062
rect 285440 144974 285620 145062
rect 285728 144974 285908 145062
rect 286016 144974 286196 145062
rect 286304 144974 286484 145062
rect 286592 144974 286772 145062
rect 286880 144974 287060 145062
rect 287314 144974 287494 145062
rect 287602 144974 287782 145062
rect 287890 144974 288070 145062
rect 288178 144974 288358 145062
rect 288466 144974 288646 145062
rect 288754 144974 288934 145062
rect 289042 144974 289222 145062
rect 289330 144974 289510 145062
rect 289764 144974 289944 145062
rect 290052 144974 290232 145062
rect 290340 144974 290520 145062
rect 290628 144974 290808 145062
rect 290916 144974 291096 145062
rect 291204 144974 291384 145062
rect 291492 144974 291672 145062
rect 291780 144974 291960 145062
rect 292214 144974 292394 145062
rect 292502 144974 292682 145062
rect 292790 144974 292970 145062
rect 293078 144974 293258 145062
rect 293366 144974 293546 145062
rect 293654 144974 293834 145062
rect 293942 144974 294122 145062
rect 294230 144974 294410 145062
rect 294664 144974 294844 145062
rect 294952 144974 295132 145062
rect 295240 144974 295420 145062
rect 295528 144974 295708 145062
rect 295816 144974 295996 145062
rect 296104 144974 296284 145062
rect 296392 144974 296572 145062
rect 296680 144974 296860 145062
rect 297114 144974 297294 145062
rect 297402 144974 297582 145062
rect 297690 144974 297870 145062
rect 297978 144974 298158 145062
rect 298266 144974 298446 145062
rect 298554 144974 298734 145062
rect 298842 144974 299022 145062
rect 299130 144974 299310 145062
rect 299564 144974 299744 145062
rect 299852 144974 300032 145062
rect 300140 144974 300320 145062
rect 300428 144974 300608 145062
rect 300716 144974 300896 145062
rect 301004 144974 301184 145062
rect 301292 144974 301472 145062
rect 301580 144974 301760 145062
rect 302014 144974 302194 145062
rect 302302 144974 302482 145062
rect 302590 144974 302770 145062
rect 302878 144974 303058 145062
rect 303166 144974 303346 145062
rect 303454 144974 303634 145062
rect 303742 144974 303922 145062
rect 304030 144974 304210 145062
rect 304464 144974 304644 145062
rect 304752 144974 304932 145062
rect 305040 144974 305220 145062
rect 305328 144974 305508 145062
rect 305616 144974 305796 145062
rect 305904 144974 306084 145062
rect 306192 144974 306372 145062
rect 306480 144974 306660 145062
rect 306914 144974 307094 145062
rect 307202 144974 307382 145062
rect 307490 144974 307670 145062
rect 307778 144974 307958 145062
rect 308066 144974 308246 145062
rect 308354 144974 308534 145062
rect 308642 144974 308822 145062
rect 308930 144974 309110 145062
rect 309364 144974 309544 145062
rect 309652 144974 309832 145062
rect 309940 144974 310120 145062
rect 310228 144974 310408 145062
rect 310516 144974 310696 145062
rect 310804 144974 310984 145062
rect 311092 144974 311272 145062
rect 311380 144974 311560 145062
rect 311814 144974 311994 145062
rect 312102 144974 312282 145062
rect 312390 144974 312570 145062
rect 312678 144974 312858 145062
rect 312966 144974 313146 145062
rect 313254 144974 313434 145062
rect 313542 144974 313722 145062
rect 313830 144974 314010 145062
rect 314264 144974 314444 145062
rect 314552 144974 314732 145062
rect 314840 144974 315020 145062
rect 315128 144974 315308 145062
rect 315416 144974 315596 145062
rect 315704 144974 315884 145062
rect 315992 144974 316172 145062
rect 316280 144974 316460 145062
rect 316714 144974 316894 145062
rect 317002 144974 317182 145062
rect 317290 144974 317470 145062
rect 317578 144974 317758 145062
rect 317866 144974 318046 145062
rect 318154 144974 318334 145062
rect 318442 144974 318622 145062
rect 318730 144974 318910 145062
rect 319164 144974 319344 145062
rect 319452 144974 319632 145062
rect 319740 144974 319920 145062
rect 320028 144974 320208 145062
rect 320316 144974 320496 145062
rect 320604 144974 320784 145062
rect 320892 144974 321072 145062
rect 321180 144974 321360 145062
rect 321614 144974 321794 145062
rect 321902 144974 322082 145062
rect 322190 144974 322370 145062
rect 322478 144974 322658 145062
rect 322766 144974 322946 145062
rect 323054 144974 323234 145062
rect 323342 144974 323522 145062
rect 323630 144974 323810 145062
rect 324064 144974 324244 145062
rect 324352 144974 324532 145062
rect 324640 144974 324820 145062
rect 324928 144974 325108 145062
rect 325216 144974 325396 145062
rect 325504 144974 325684 145062
rect 325792 144974 325972 145062
rect 326080 144974 326260 145062
rect 326514 144974 326694 145062
rect 326802 144974 326982 145062
rect 327090 144974 327270 145062
rect 327378 144974 327558 145062
rect 327666 144974 327846 145062
rect 327954 144974 328134 145062
rect 328242 144974 328422 145062
rect 328530 144974 328710 145062
rect 328964 144974 329144 145062
rect 329252 144974 329432 145062
rect 329540 144974 329720 145062
rect 329828 144974 330008 145062
rect 330116 144974 330296 145062
rect 330404 144974 330584 145062
rect 330692 144974 330872 145062
rect 330980 144974 331160 145062
rect 331414 144974 331594 145062
rect 331702 144974 331882 145062
rect 331990 144974 332170 145062
rect 332278 144974 332458 145062
rect 332566 144974 332746 145062
rect 332854 144974 333034 145062
rect 333142 144974 333322 145062
rect 333430 144974 333610 145062
rect 333864 144974 334044 145062
rect 334152 144974 334332 145062
rect 334440 144974 334620 145062
rect 334728 144974 334908 145062
rect 335016 144974 335196 145062
rect 335304 144974 335484 145062
rect 335592 144974 335772 145062
rect 335880 144974 336060 145062
rect 336314 144974 336494 145062
rect 336602 144974 336782 145062
rect 336890 144974 337070 145062
rect 337178 144974 337358 145062
rect 337466 144974 337646 145062
rect 337754 144974 337934 145062
rect 338042 144974 338222 145062
rect 338330 144974 338510 145062
rect 338764 144974 338944 145062
rect 339052 144974 339232 145062
rect 339340 144974 339520 145062
rect 339628 144974 339808 145062
rect 339916 144974 340096 145062
rect 340204 144974 340384 145062
rect 340492 144974 340672 145062
rect 340780 144974 340960 145062
rect 341214 144974 341394 145062
rect 341502 144974 341682 145062
rect 341790 144974 341970 145062
rect 342078 144974 342258 145062
rect 342366 144974 342546 145062
rect 342654 144974 342834 145062
rect 342942 144974 343122 145062
rect 343230 144974 343410 145062
rect 343664 144974 343844 145062
rect 343952 144974 344132 145062
rect 344240 144974 344420 145062
rect 344528 144974 344708 145062
rect 344816 144974 344996 145062
rect 345104 144974 345284 145062
rect 345392 144974 345572 145062
rect 345680 144974 345860 145062
rect 346114 144974 346294 145062
rect 346402 144974 346582 145062
rect 346690 144974 346870 145062
rect 346978 144974 347158 145062
rect 347266 144974 347446 145062
rect 347554 144974 347734 145062
rect 347842 144974 348022 145062
rect 348130 144974 348310 145062
rect 348564 144974 348744 145062
rect 348852 144974 349032 145062
rect 349140 144974 349320 145062
rect 349428 144974 349608 145062
rect 349716 144974 349896 145062
rect 350004 144974 350184 145062
rect 350292 144974 350472 145062
rect 350580 144974 350760 145062
rect 351014 144974 351194 145062
rect 351302 144974 351482 145062
rect 351590 144974 351770 145062
rect 351878 144974 352058 145062
rect 352166 144974 352346 145062
rect 352454 144974 352634 145062
rect 352742 144974 352922 145062
rect 353030 144974 353210 145062
rect 353464 144974 353644 145062
rect 353752 144974 353932 145062
rect 354040 144974 354220 145062
rect 354328 144974 354508 145062
rect 354616 144974 354796 145062
rect 354904 144974 355084 145062
rect 355192 144974 355372 145062
rect 355480 144974 355660 145062
rect 355914 144974 356094 145062
rect 356202 144974 356382 145062
rect 356490 144974 356670 145062
rect 356778 144974 356958 145062
rect 357066 144974 357246 145062
rect 357354 144974 357534 145062
rect 357642 144974 357822 145062
rect 357930 144974 358110 145062
rect 358364 144974 358544 145062
rect 358652 144974 358832 145062
rect 358940 144974 359120 145062
rect 359228 144974 359408 145062
rect 359516 144974 359696 145062
rect 359804 144974 359984 145062
rect 360092 144974 360272 145062
rect 360380 144974 360560 145062
rect 360814 144974 360994 145062
rect 361102 144974 361282 145062
rect 361390 144974 361570 145062
rect 361678 144974 361858 145062
rect 361966 144974 362146 145062
rect 362254 144974 362434 145062
rect 362542 144974 362722 145062
rect 362830 144974 363010 145062
rect 363264 144974 363444 145062
rect 363552 144974 363732 145062
rect 363840 144974 364020 145062
rect 364128 144974 364308 145062
rect 364416 144974 364596 145062
rect 364704 144974 364884 145062
rect 364992 144974 365172 145062
rect 365280 144974 365460 145062
rect 365714 144974 365894 145062
rect 366002 144974 366182 145062
rect 366290 144974 366470 145062
rect 366578 144974 366758 145062
rect 366866 144974 367046 145062
rect 367154 144974 367334 145062
rect 367442 144974 367622 145062
rect 367730 144974 367910 145062
rect 243214 144758 243394 144846
rect 243502 144758 243682 144846
rect 243790 144758 243970 144846
rect 244078 144758 244258 144846
rect 244366 144758 244546 144846
rect 244654 144758 244834 144846
rect 244942 144758 245122 144846
rect 245230 144758 245410 144846
rect 245664 144758 245844 144846
rect 245952 144758 246132 144846
rect 246240 144758 246420 144846
rect 246528 144758 246708 144846
rect 246816 144758 246996 144846
rect 247104 144758 247284 144846
rect 247392 144758 247572 144846
rect 247680 144758 247860 144846
rect 248114 144758 248294 144846
rect 248402 144758 248582 144846
rect 248690 144758 248870 144846
rect 248978 144758 249158 144846
rect 249266 144758 249446 144846
rect 249554 144758 249734 144846
rect 249842 144758 250022 144846
rect 250130 144758 250310 144846
rect 250564 144758 250744 144846
rect 250852 144758 251032 144846
rect 251140 144758 251320 144846
rect 251428 144758 251608 144846
rect 251716 144758 251896 144846
rect 252004 144758 252184 144846
rect 252292 144758 252472 144846
rect 252580 144758 252760 144846
rect 253014 144758 253194 144846
rect 253302 144758 253482 144846
rect 253590 144758 253770 144846
rect 253878 144758 254058 144846
rect 254166 144758 254346 144846
rect 254454 144758 254634 144846
rect 254742 144758 254922 144846
rect 255030 144758 255210 144846
rect 255464 144758 255644 144846
rect 255752 144758 255932 144846
rect 256040 144758 256220 144846
rect 256328 144758 256508 144846
rect 256616 144758 256796 144846
rect 256904 144758 257084 144846
rect 257192 144758 257372 144846
rect 257480 144758 257660 144846
rect 257914 144758 258094 144846
rect 258202 144758 258382 144846
rect 258490 144758 258670 144846
rect 258778 144758 258958 144846
rect 259066 144758 259246 144846
rect 259354 144758 259534 144846
rect 259642 144758 259822 144846
rect 259930 144758 260110 144846
rect 260364 144758 260544 144846
rect 260652 144758 260832 144846
rect 260940 144758 261120 144846
rect 261228 144758 261408 144846
rect 261516 144758 261696 144846
rect 261804 144758 261984 144846
rect 262092 144758 262272 144846
rect 262380 144758 262560 144846
rect 262814 144758 262994 144846
rect 263102 144758 263282 144846
rect 263390 144758 263570 144846
rect 263678 144758 263858 144846
rect 263966 144758 264146 144846
rect 264254 144758 264434 144846
rect 264542 144758 264722 144846
rect 264830 144758 265010 144846
rect 265264 144758 265444 144846
rect 265552 144758 265732 144846
rect 265840 144758 266020 144846
rect 266128 144758 266308 144846
rect 266416 144758 266596 144846
rect 266704 144758 266884 144846
rect 266992 144758 267172 144846
rect 267280 144758 267460 144846
rect 267714 144758 267894 144846
rect 268002 144758 268182 144846
rect 268290 144758 268470 144846
rect 268578 144758 268758 144846
rect 268866 144758 269046 144846
rect 269154 144758 269334 144846
rect 269442 144758 269622 144846
rect 269730 144758 269910 144846
rect 270164 144758 270344 144846
rect 270452 144758 270632 144846
rect 270740 144758 270920 144846
rect 271028 144758 271208 144846
rect 271316 144758 271496 144846
rect 271604 144758 271784 144846
rect 271892 144758 272072 144846
rect 272180 144758 272360 144846
rect 272614 144758 272794 144846
rect 272902 144758 273082 144846
rect 273190 144758 273370 144846
rect 273478 144758 273658 144846
rect 273766 144758 273946 144846
rect 274054 144758 274234 144846
rect 274342 144758 274522 144846
rect 274630 144758 274810 144846
rect 275064 144758 275244 144846
rect 275352 144758 275532 144846
rect 275640 144758 275820 144846
rect 275928 144758 276108 144846
rect 276216 144758 276396 144846
rect 276504 144758 276684 144846
rect 276792 144758 276972 144846
rect 277080 144758 277260 144846
rect 277514 144758 277694 144846
rect 277802 144758 277982 144846
rect 278090 144758 278270 144846
rect 278378 144758 278558 144846
rect 278666 144758 278846 144846
rect 278954 144758 279134 144846
rect 279242 144758 279422 144846
rect 279530 144758 279710 144846
rect 279964 144758 280144 144846
rect 280252 144758 280432 144846
rect 280540 144758 280720 144846
rect 280828 144758 281008 144846
rect 281116 144758 281296 144846
rect 281404 144758 281584 144846
rect 281692 144758 281872 144846
rect 281980 144758 282160 144846
rect 282414 144758 282594 144846
rect 282702 144758 282882 144846
rect 282990 144758 283170 144846
rect 283278 144758 283458 144846
rect 283566 144758 283746 144846
rect 283854 144758 284034 144846
rect 284142 144758 284322 144846
rect 284430 144758 284610 144846
rect 284864 144758 285044 144846
rect 285152 144758 285332 144846
rect 285440 144758 285620 144846
rect 285728 144758 285908 144846
rect 286016 144758 286196 144846
rect 286304 144758 286484 144846
rect 286592 144758 286772 144846
rect 286880 144758 287060 144846
rect 287314 144758 287494 144846
rect 287602 144758 287782 144846
rect 287890 144758 288070 144846
rect 288178 144758 288358 144846
rect 288466 144758 288646 144846
rect 288754 144758 288934 144846
rect 289042 144758 289222 144846
rect 289330 144758 289510 144846
rect 289764 144758 289944 144846
rect 290052 144758 290232 144846
rect 290340 144758 290520 144846
rect 290628 144758 290808 144846
rect 290916 144758 291096 144846
rect 291204 144758 291384 144846
rect 291492 144758 291672 144846
rect 291780 144758 291960 144846
rect 292214 144758 292394 144846
rect 292502 144758 292682 144846
rect 292790 144758 292970 144846
rect 293078 144758 293258 144846
rect 293366 144758 293546 144846
rect 293654 144758 293834 144846
rect 293942 144758 294122 144846
rect 294230 144758 294410 144846
rect 294664 144758 294844 144846
rect 294952 144758 295132 144846
rect 295240 144758 295420 144846
rect 295528 144758 295708 144846
rect 295816 144758 295996 144846
rect 296104 144758 296284 144846
rect 296392 144758 296572 144846
rect 296680 144758 296860 144846
rect 297114 144758 297294 144846
rect 297402 144758 297582 144846
rect 297690 144758 297870 144846
rect 297978 144758 298158 144846
rect 298266 144758 298446 144846
rect 298554 144758 298734 144846
rect 298842 144758 299022 144846
rect 299130 144758 299310 144846
rect 299564 144758 299744 144846
rect 299852 144758 300032 144846
rect 300140 144758 300320 144846
rect 300428 144758 300608 144846
rect 300716 144758 300896 144846
rect 301004 144758 301184 144846
rect 301292 144758 301472 144846
rect 301580 144758 301760 144846
rect 302014 144758 302194 144846
rect 302302 144758 302482 144846
rect 302590 144758 302770 144846
rect 302878 144758 303058 144846
rect 303166 144758 303346 144846
rect 303454 144758 303634 144846
rect 303742 144758 303922 144846
rect 304030 144758 304210 144846
rect 304464 144758 304644 144846
rect 304752 144758 304932 144846
rect 305040 144758 305220 144846
rect 305328 144758 305508 144846
rect 305616 144758 305796 144846
rect 305904 144758 306084 144846
rect 306192 144758 306372 144846
rect 306480 144758 306660 144846
rect 306914 144758 307094 144846
rect 307202 144758 307382 144846
rect 307490 144758 307670 144846
rect 307778 144758 307958 144846
rect 308066 144758 308246 144846
rect 308354 144758 308534 144846
rect 308642 144758 308822 144846
rect 308930 144758 309110 144846
rect 309364 144758 309544 144846
rect 309652 144758 309832 144846
rect 309940 144758 310120 144846
rect 310228 144758 310408 144846
rect 310516 144758 310696 144846
rect 310804 144758 310984 144846
rect 311092 144758 311272 144846
rect 311380 144758 311560 144846
rect 311814 144758 311994 144846
rect 312102 144758 312282 144846
rect 312390 144758 312570 144846
rect 312678 144758 312858 144846
rect 312966 144758 313146 144846
rect 313254 144758 313434 144846
rect 313542 144758 313722 144846
rect 313830 144758 314010 144846
rect 314264 144758 314444 144846
rect 314552 144758 314732 144846
rect 314840 144758 315020 144846
rect 315128 144758 315308 144846
rect 315416 144758 315596 144846
rect 315704 144758 315884 144846
rect 315992 144758 316172 144846
rect 316280 144758 316460 144846
rect 316714 144758 316894 144846
rect 317002 144758 317182 144846
rect 317290 144758 317470 144846
rect 317578 144758 317758 144846
rect 317866 144758 318046 144846
rect 318154 144758 318334 144846
rect 318442 144758 318622 144846
rect 318730 144758 318910 144846
rect 319164 144758 319344 144846
rect 319452 144758 319632 144846
rect 319740 144758 319920 144846
rect 320028 144758 320208 144846
rect 320316 144758 320496 144846
rect 320604 144758 320784 144846
rect 320892 144758 321072 144846
rect 321180 144758 321360 144846
rect 321614 144758 321794 144846
rect 321902 144758 322082 144846
rect 322190 144758 322370 144846
rect 322478 144758 322658 144846
rect 322766 144758 322946 144846
rect 323054 144758 323234 144846
rect 323342 144758 323522 144846
rect 323630 144758 323810 144846
rect 324064 144758 324244 144846
rect 324352 144758 324532 144846
rect 324640 144758 324820 144846
rect 324928 144758 325108 144846
rect 325216 144758 325396 144846
rect 325504 144758 325684 144846
rect 325792 144758 325972 144846
rect 326080 144758 326260 144846
rect 326514 144758 326694 144846
rect 326802 144758 326982 144846
rect 327090 144758 327270 144846
rect 327378 144758 327558 144846
rect 327666 144758 327846 144846
rect 327954 144758 328134 144846
rect 328242 144758 328422 144846
rect 328530 144758 328710 144846
rect 328964 144758 329144 144846
rect 329252 144758 329432 144846
rect 329540 144758 329720 144846
rect 329828 144758 330008 144846
rect 330116 144758 330296 144846
rect 330404 144758 330584 144846
rect 330692 144758 330872 144846
rect 330980 144758 331160 144846
rect 331414 144758 331594 144846
rect 331702 144758 331882 144846
rect 331990 144758 332170 144846
rect 332278 144758 332458 144846
rect 332566 144758 332746 144846
rect 332854 144758 333034 144846
rect 333142 144758 333322 144846
rect 333430 144758 333610 144846
rect 333864 144758 334044 144846
rect 334152 144758 334332 144846
rect 334440 144758 334620 144846
rect 334728 144758 334908 144846
rect 335016 144758 335196 144846
rect 335304 144758 335484 144846
rect 335592 144758 335772 144846
rect 335880 144758 336060 144846
rect 336314 144758 336494 144846
rect 336602 144758 336782 144846
rect 336890 144758 337070 144846
rect 337178 144758 337358 144846
rect 337466 144758 337646 144846
rect 337754 144758 337934 144846
rect 338042 144758 338222 144846
rect 338330 144758 338510 144846
rect 338764 144758 338944 144846
rect 339052 144758 339232 144846
rect 339340 144758 339520 144846
rect 339628 144758 339808 144846
rect 339916 144758 340096 144846
rect 340204 144758 340384 144846
rect 340492 144758 340672 144846
rect 340780 144758 340960 144846
rect 341214 144758 341394 144846
rect 341502 144758 341682 144846
rect 341790 144758 341970 144846
rect 342078 144758 342258 144846
rect 342366 144758 342546 144846
rect 342654 144758 342834 144846
rect 342942 144758 343122 144846
rect 343230 144758 343410 144846
rect 343664 144758 343844 144846
rect 343952 144758 344132 144846
rect 344240 144758 344420 144846
rect 344528 144758 344708 144846
rect 344816 144758 344996 144846
rect 345104 144758 345284 144846
rect 345392 144758 345572 144846
rect 345680 144758 345860 144846
rect 346114 144758 346294 144846
rect 346402 144758 346582 144846
rect 346690 144758 346870 144846
rect 346978 144758 347158 144846
rect 347266 144758 347446 144846
rect 347554 144758 347734 144846
rect 347842 144758 348022 144846
rect 348130 144758 348310 144846
rect 348564 144758 348744 144846
rect 348852 144758 349032 144846
rect 349140 144758 349320 144846
rect 349428 144758 349608 144846
rect 349716 144758 349896 144846
rect 350004 144758 350184 144846
rect 350292 144758 350472 144846
rect 350580 144758 350760 144846
rect 351014 144758 351194 144846
rect 351302 144758 351482 144846
rect 351590 144758 351770 144846
rect 351878 144758 352058 144846
rect 352166 144758 352346 144846
rect 352454 144758 352634 144846
rect 352742 144758 352922 144846
rect 353030 144758 353210 144846
rect 353464 144758 353644 144846
rect 353752 144758 353932 144846
rect 354040 144758 354220 144846
rect 354328 144758 354508 144846
rect 354616 144758 354796 144846
rect 354904 144758 355084 144846
rect 355192 144758 355372 144846
rect 355480 144758 355660 144846
rect 355914 144758 356094 144846
rect 356202 144758 356382 144846
rect 356490 144758 356670 144846
rect 356778 144758 356958 144846
rect 357066 144758 357246 144846
rect 357354 144758 357534 144846
rect 357642 144758 357822 144846
rect 357930 144758 358110 144846
rect 358364 144758 358544 144846
rect 358652 144758 358832 144846
rect 358940 144758 359120 144846
rect 359228 144758 359408 144846
rect 359516 144758 359696 144846
rect 359804 144758 359984 144846
rect 360092 144758 360272 144846
rect 360380 144758 360560 144846
rect 360814 144758 360994 144846
rect 361102 144758 361282 144846
rect 361390 144758 361570 144846
rect 361678 144758 361858 144846
rect 361966 144758 362146 144846
rect 362254 144758 362434 144846
rect 362542 144758 362722 144846
rect 362830 144758 363010 144846
rect 363264 144758 363444 144846
rect 363552 144758 363732 144846
rect 363840 144758 364020 144846
rect 364128 144758 364308 144846
rect 364416 144758 364596 144846
rect 364704 144758 364884 144846
rect 364992 144758 365172 144846
rect 365280 144758 365460 144846
rect 365714 144758 365894 144846
rect 366002 144758 366182 144846
rect 366290 144758 366470 144846
rect 366578 144758 366758 144846
rect 366866 144758 367046 144846
rect 367154 144758 367334 144846
rect 367442 144758 367622 144846
rect 367730 144758 367910 144846
rect 243214 144282 243394 144370
rect 243502 144282 243682 144370
rect 243790 144282 243970 144370
rect 244078 144282 244258 144370
rect 244366 144282 244546 144370
rect 244654 144282 244834 144370
rect 244942 144282 245122 144370
rect 245230 144282 245410 144370
rect 245664 144282 245844 144370
rect 245952 144282 246132 144370
rect 246240 144282 246420 144370
rect 246528 144282 246708 144370
rect 246816 144282 246996 144370
rect 247104 144282 247284 144370
rect 247392 144282 247572 144370
rect 247680 144282 247860 144370
rect 248114 144282 248294 144370
rect 248402 144282 248582 144370
rect 248690 144282 248870 144370
rect 248978 144282 249158 144370
rect 249266 144282 249446 144370
rect 249554 144282 249734 144370
rect 249842 144282 250022 144370
rect 250130 144282 250310 144370
rect 250564 144282 250744 144370
rect 250852 144282 251032 144370
rect 251140 144282 251320 144370
rect 251428 144282 251608 144370
rect 251716 144282 251896 144370
rect 252004 144282 252184 144370
rect 252292 144282 252472 144370
rect 252580 144282 252760 144370
rect 253014 144282 253194 144370
rect 253302 144282 253482 144370
rect 253590 144282 253770 144370
rect 253878 144282 254058 144370
rect 254166 144282 254346 144370
rect 254454 144282 254634 144370
rect 254742 144282 254922 144370
rect 255030 144282 255210 144370
rect 255464 144282 255644 144370
rect 255752 144282 255932 144370
rect 256040 144282 256220 144370
rect 256328 144282 256508 144370
rect 256616 144282 256796 144370
rect 256904 144282 257084 144370
rect 257192 144282 257372 144370
rect 257480 144282 257660 144370
rect 257914 144282 258094 144370
rect 258202 144282 258382 144370
rect 258490 144282 258670 144370
rect 258778 144282 258958 144370
rect 259066 144282 259246 144370
rect 259354 144282 259534 144370
rect 259642 144282 259822 144370
rect 259930 144282 260110 144370
rect 260364 144282 260544 144370
rect 260652 144282 260832 144370
rect 260940 144282 261120 144370
rect 261228 144282 261408 144370
rect 261516 144282 261696 144370
rect 261804 144282 261984 144370
rect 262092 144282 262272 144370
rect 262380 144282 262560 144370
rect 262814 144282 262994 144370
rect 263102 144282 263282 144370
rect 263390 144282 263570 144370
rect 263678 144282 263858 144370
rect 263966 144282 264146 144370
rect 264254 144282 264434 144370
rect 264542 144282 264722 144370
rect 264830 144282 265010 144370
rect 265264 144282 265444 144370
rect 265552 144282 265732 144370
rect 265840 144282 266020 144370
rect 266128 144282 266308 144370
rect 266416 144282 266596 144370
rect 266704 144282 266884 144370
rect 266992 144282 267172 144370
rect 267280 144282 267460 144370
rect 267714 144282 267894 144370
rect 268002 144282 268182 144370
rect 268290 144282 268470 144370
rect 268578 144282 268758 144370
rect 268866 144282 269046 144370
rect 269154 144282 269334 144370
rect 269442 144282 269622 144370
rect 269730 144282 269910 144370
rect 270164 144282 270344 144370
rect 270452 144282 270632 144370
rect 270740 144282 270920 144370
rect 271028 144282 271208 144370
rect 271316 144282 271496 144370
rect 271604 144282 271784 144370
rect 271892 144282 272072 144370
rect 272180 144282 272360 144370
rect 272614 144282 272794 144370
rect 272902 144282 273082 144370
rect 273190 144282 273370 144370
rect 273478 144282 273658 144370
rect 273766 144282 273946 144370
rect 274054 144282 274234 144370
rect 274342 144282 274522 144370
rect 274630 144282 274810 144370
rect 275064 144282 275244 144370
rect 275352 144282 275532 144370
rect 275640 144282 275820 144370
rect 275928 144282 276108 144370
rect 276216 144282 276396 144370
rect 276504 144282 276684 144370
rect 276792 144282 276972 144370
rect 277080 144282 277260 144370
rect 277514 144282 277694 144370
rect 277802 144282 277982 144370
rect 278090 144282 278270 144370
rect 278378 144282 278558 144370
rect 278666 144282 278846 144370
rect 278954 144282 279134 144370
rect 279242 144282 279422 144370
rect 279530 144282 279710 144370
rect 279964 144282 280144 144370
rect 280252 144282 280432 144370
rect 280540 144282 280720 144370
rect 280828 144282 281008 144370
rect 281116 144282 281296 144370
rect 281404 144282 281584 144370
rect 281692 144282 281872 144370
rect 281980 144282 282160 144370
rect 282414 144282 282594 144370
rect 282702 144282 282882 144370
rect 282990 144282 283170 144370
rect 283278 144282 283458 144370
rect 283566 144282 283746 144370
rect 283854 144282 284034 144370
rect 284142 144282 284322 144370
rect 284430 144282 284610 144370
rect 284864 144282 285044 144370
rect 285152 144282 285332 144370
rect 285440 144282 285620 144370
rect 285728 144282 285908 144370
rect 286016 144282 286196 144370
rect 286304 144282 286484 144370
rect 286592 144282 286772 144370
rect 286880 144282 287060 144370
rect 287314 144282 287494 144370
rect 287602 144282 287782 144370
rect 287890 144282 288070 144370
rect 288178 144282 288358 144370
rect 288466 144282 288646 144370
rect 288754 144282 288934 144370
rect 289042 144282 289222 144370
rect 289330 144282 289510 144370
rect 289764 144282 289944 144370
rect 290052 144282 290232 144370
rect 290340 144282 290520 144370
rect 290628 144282 290808 144370
rect 290916 144282 291096 144370
rect 291204 144282 291384 144370
rect 291492 144282 291672 144370
rect 291780 144282 291960 144370
rect 292214 144282 292394 144370
rect 292502 144282 292682 144370
rect 292790 144282 292970 144370
rect 293078 144282 293258 144370
rect 293366 144282 293546 144370
rect 293654 144282 293834 144370
rect 293942 144282 294122 144370
rect 294230 144282 294410 144370
rect 294664 144282 294844 144370
rect 294952 144282 295132 144370
rect 295240 144282 295420 144370
rect 295528 144282 295708 144370
rect 295816 144282 295996 144370
rect 296104 144282 296284 144370
rect 296392 144282 296572 144370
rect 296680 144282 296860 144370
rect 297114 144282 297294 144370
rect 297402 144282 297582 144370
rect 297690 144282 297870 144370
rect 297978 144282 298158 144370
rect 298266 144282 298446 144370
rect 298554 144282 298734 144370
rect 298842 144282 299022 144370
rect 299130 144282 299310 144370
rect 299564 144282 299744 144370
rect 299852 144282 300032 144370
rect 300140 144282 300320 144370
rect 300428 144282 300608 144370
rect 300716 144282 300896 144370
rect 301004 144282 301184 144370
rect 301292 144282 301472 144370
rect 301580 144282 301760 144370
rect 302014 144282 302194 144370
rect 302302 144282 302482 144370
rect 302590 144282 302770 144370
rect 302878 144282 303058 144370
rect 303166 144282 303346 144370
rect 303454 144282 303634 144370
rect 303742 144282 303922 144370
rect 304030 144282 304210 144370
rect 304464 144282 304644 144370
rect 304752 144282 304932 144370
rect 305040 144282 305220 144370
rect 305328 144282 305508 144370
rect 305616 144282 305796 144370
rect 305904 144282 306084 144370
rect 306192 144282 306372 144370
rect 306480 144282 306660 144370
rect 306914 144282 307094 144370
rect 307202 144282 307382 144370
rect 307490 144282 307670 144370
rect 307778 144282 307958 144370
rect 308066 144282 308246 144370
rect 308354 144282 308534 144370
rect 308642 144282 308822 144370
rect 308930 144282 309110 144370
rect 309364 144282 309544 144370
rect 309652 144282 309832 144370
rect 309940 144282 310120 144370
rect 310228 144282 310408 144370
rect 310516 144282 310696 144370
rect 310804 144282 310984 144370
rect 311092 144282 311272 144370
rect 311380 144282 311560 144370
rect 311814 144282 311994 144370
rect 312102 144282 312282 144370
rect 312390 144282 312570 144370
rect 312678 144282 312858 144370
rect 312966 144282 313146 144370
rect 313254 144282 313434 144370
rect 313542 144282 313722 144370
rect 313830 144282 314010 144370
rect 314264 144282 314444 144370
rect 314552 144282 314732 144370
rect 314840 144282 315020 144370
rect 315128 144282 315308 144370
rect 315416 144282 315596 144370
rect 315704 144282 315884 144370
rect 315992 144282 316172 144370
rect 316280 144282 316460 144370
rect 316714 144282 316894 144370
rect 317002 144282 317182 144370
rect 317290 144282 317470 144370
rect 317578 144282 317758 144370
rect 317866 144282 318046 144370
rect 318154 144282 318334 144370
rect 318442 144282 318622 144370
rect 318730 144282 318910 144370
rect 319164 144282 319344 144370
rect 319452 144282 319632 144370
rect 319740 144282 319920 144370
rect 320028 144282 320208 144370
rect 320316 144282 320496 144370
rect 320604 144282 320784 144370
rect 320892 144282 321072 144370
rect 321180 144282 321360 144370
rect 321614 144282 321794 144370
rect 321902 144282 322082 144370
rect 322190 144282 322370 144370
rect 322478 144282 322658 144370
rect 322766 144282 322946 144370
rect 323054 144282 323234 144370
rect 323342 144282 323522 144370
rect 323630 144282 323810 144370
rect 324064 144282 324244 144370
rect 324352 144282 324532 144370
rect 324640 144282 324820 144370
rect 324928 144282 325108 144370
rect 325216 144282 325396 144370
rect 325504 144282 325684 144370
rect 325792 144282 325972 144370
rect 326080 144282 326260 144370
rect 326514 144282 326694 144370
rect 326802 144282 326982 144370
rect 327090 144282 327270 144370
rect 327378 144282 327558 144370
rect 327666 144282 327846 144370
rect 327954 144282 328134 144370
rect 328242 144282 328422 144370
rect 328530 144282 328710 144370
rect 328964 144282 329144 144370
rect 329252 144282 329432 144370
rect 329540 144282 329720 144370
rect 329828 144282 330008 144370
rect 330116 144282 330296 144370
rect 330404 144282 330584 144370
rect 330692 144282 330872 144370
rect 330980 144282 331160 144370
rect 331414 144282 331594 144370
rect 331702 144282 331882 144370
rect 331990 144282 332170 144370
rect 332278 144282 332458 144370
rect 332566 144282 332746 144370
rect 332854 144282 333034 144370
rect 333142 144282 333322 144370
rect 333430 144282 333610 144370
rect 333864 144282 334044 144370
rect 334152 144282 334332 144370
rect 334440 144282 334620 144370
rect 334728 144282 334908 144370
rect 335016 144282 335196 144370
rect 335304 144282 335484 144370
rect 335592 144282 335772 144370
rect 335880 144282 336060 144370
rect 336314 144282 336494 144370
rect 336602 144282 336782 144370
rect 336890 144282 337070 144370
rect 337178 144282 337358 144370
rect 337466 144282 337646 144370
rect 337754 144282 337934 144370
rect 338042 144282 338222 144370
rect 338330 144282 338510 144370
rect 338764 144282 338944 144370
rect 339052 144282 339232 144370
rect 339340 144282 339520 144370
rect 339628 144282 339808 144370
rect 339916 144282 340096 144370
rect 340204 144282 340384 144370
rect 340492 144282 340672 144370
rect 340780 144282 340960 144370
rect 341214 144282 341394 144370
rect 341502 144282 341682 144370
rect 341790 144282 341970 144370
rect 342078 144282 342258 144370
rect 342366 144282 342546 144370
rect 342654 144282 342834 144370
rect 342942 144282 343122 144370
rect 343230 144282 343410 144370
rect 343664 144282 343844 144370
rect 343952 144282 344132 144370
rect 344240 144282 344420 144370
rect 344528 144282 344708 144370
rect 344816 144282 344996 144370
rect 345104 144282 345284 144370
rect 345392 144282 345572 144370
rect 345680 144282 345860 144370
rect 346114 144282 346294 144370
rect 346402 144282 346582 144370
rect 346690 144282 346870 144370
rect 346978 144282 347158 144370
rect 347266 144282 347446 144370
rect 347554 144282 347734 144370
rect 347842 144282 348022 144370
rect 348130 144282 348310 144370
rect 348564 144282 348744 144370
rect 348852 144282 349032 144370
rect 349140 144282 349320 144370
rect 349428 144282 349608 144370
rect 349716 144282 349896 144370
rect 350004 144282 350184 144370
rect 350292 144282 350472 144370
rect 350580 144282 350760 144370
rect 351014 144282 351194 144370
rect 351302 144282 351482 144370
rect 351590 144282 351770 144370
rect 351878 144282 352058 144370
rect 352166 144282 352346 144370
rect 352454 144282 352634 144370
rect 352742 144282 352922 144370
rect 353030 144282 353210 144370
rect 353464 144282 353644 144370
rect 353752 144282 353932 144370
rect 354040 144282 354220 144370
rect 354328 144282 354508 144370
rect 354616 144282 354796 144370
rect 354904 144282 355084 144370
rect 355192 144282 355372 144370
rect 355480 144282 355660 144370
rect 355914 144282 356094 144370
rect 356202 144282 356382 144370
rect 356490 144282 356670 144370
rect 356778 144282 356958 144370
rect 357066 144282 357246 144370
rect 357354 144282 357534 144370
rect 357642 144282 357822 144370
rect 357930 144282 358110 144370
rect 358364 144282 358544 144370
rect 358652 144282 358832 144370
rect 358940 144282 359120 144370
rect 359228 144282 359408 144370
rect 359516 144282 359696 144370
rect 359804 144282 359984 144370
rect 360092 144282 360272 144370
rect 360380 144282 360560 144370
rect 360814 144282 360994 144370
rect 361102 144282 361282 144370
rect 361390 144282 361570 144370
rect 361678 144282 361858 144370
rect 361966 144282 362146 144370
rect 362254 144282 362434 144370
rect 362542 144282 362722 144370
rect 362830 144282 363010 144370
rect 363264 144282 363444 144370
rect 363552 144282 363732 144370
rect 363840 144282 364020 144370
rect 364128 144282 364308 144370
rect 364416 144282 364596 144370
rect 364704 144282 364884 144370
rect 364992 144282 365172 144370
rect 365280 144282 365460 144370
rect 365714 144282 365894 144370
rect 366002 144282 366182 144370
rect 366290 144282 366470 144370
rect 366578 144282 366758 144370
rect 366866 144282 367046 144370
rect 367154 144282 367334 144370
rect 367442 144282 367622 144370
rect 367730 144282 367910 144370
rect 243214 144066 243394 144154
rect 243502 144066 243682 144154
rect 243790 144066 243970 144154
rect 244078 144066 244258 144154
rect 244366 144066 244546 144154
rect 244654 144066 244834 144154
rect 244942 144066 245122 144154
rect 245230 144066 245410 144154
rect 245664 144066 245844 144154
rect 245952 144066 246132 144154
rect 246240 144066 246420 144154
rect 246528 144066 246708 144154
rect 246816 144066 246996 144154
rect 247104 144066 247284 144154
rect 247392 144066 247572 144154
rect 247680 144066 247860 144154
rect 248114 144066 248294 144154
rect 248402 144066 248582 144154
rect 248690 144066 248870 144154
rect 248978 144066 249158 144154
rect 249266 144066 249446 144154
rect 249554 144066 249734 144154
rect 249842 144066 250022 144154
rect 250130 144066 250310 144154
rect 250564 144066 250744 144154
rect 250852 144066 251032 144154
rect 251140 144066 251320 144154
rect 251428 144066 251608 144154
rect 251716 144066 251896 144154
rect 252004 144066 252184 144154
rect 252292 144066 252472 144154
rect 252580 144066 252760 144154
rect 253014 144066 253194 144154
rect 253302 144066 253482 144154
rect 253590 144066 253770 144154
rect 253878 144066 254058 144154
rect 254166 144066 254346 144154
rect 254454 144066 254634 144154
rect 254742 144066 254922 144154
rect 255030 144066 255210 144154
rect 255464 144066 255644 144154
rect 255752 144066 255932 144154
rect 256040 144066 256220 144154
rect 256328 144066 256508 144154
rect 256616 144066 256796 144154
rect 256904 144066 257084 144154
rect 257192 144066 257372 144154
rect 257480 144066 257660 144154
rect 257914 144066 258094 144154
rect 258202 144066 258382 144154
rect 258490 144066 258670 144154
rect 258778 144066 258958 144154
rect 259066 144066 259246 144154
rect 259354 144066 259534 144154
rect 259642 144066 259822 144154
rect 259930 144066 260110 144154
rect 260364 144066 260544 144154
rect 260652 144066 260832 144154
rect 260940 144066 261120 144154
rect 261228 144066 261408 144154
rect 261516 144066 261696 144154
rect 261804 144066 261984 144154
rect 262092 144066 262272 144154
rect 262380 144066 262560 144154
rect 262814 144066 262994 144154
rect 263102 144066 263282 144154
rect 263390 144066 263570 144154
rect 263678 144066 263858 144154
rect 263966 144066 264146 144154
rect 264254 144066 264434 144154
rect 264542 144066 264722 144154
rect 264830 144066 265010 144154
rect 265264 144066 265444 144154
rect 265552 144066 265732 144154
rect 265840 144066 266020 144154
rect 266128 144066 266308 144154
rect 266416 144066 266596 144154
rect 266704 144066 266884 144154
rect 266992 144066 267172 144154
rect 267280 144066 267460 144154
rect 267714 144066 267894 144154
rect 268002 144066 268182 144154
rect 268290 144066 268470 144154
rect 268578 144066 268758 144154
rect 268866 144066 269046 144154
rect 269154 144066 269334 144154
rect 269442 144066 269622 144154
rect 269730 144066 269910 144154
rect 270164 144066 270344 144154
rect 270452 144066 270632 144154
rect 270740 144066 270920 144154
rect 271028 144066 271208 144154
rect 271316 144066 271496 144154
rect 271604 144066 271784 144154
rect 271892 144066 272072 144154
rect 272180 144066 272360 144154
rect 272614 144066 272794 144154
rect 272902 144066 273082 144154
rect 273190 144066 273370 144154
rect 273478 144066 273658 144154
rect 273766 144066 273946 144154
rect 274054 144066 274234 144154
rect 274342 144066 274522 144154
rect 274630 144066 274810 144154
rect 275064 144066 275244 144154
rect 275352 144066 275532 144154
rect 275640 144066 275820 144154
rect 275928 144066 276108 144154
rect 276216 144066 276396 144154
rect 276504 144066 276684 144154
rect 276792 144066 276972 144154
rect 277080 144066 277260 144154
rect 277514 144066 277694 144154
rect 277802 144066 277982 144154
rect 278090 144066 278270 144154
rect 278378 144066 278558 144154
rect 278666 144066 278846 144154
rect 278954 144066 279134 144154
rect 279242 144066 279422 144154
rect 279530 144066 279710 144154
rect 279964 144066 280144 144154
rect 280252 144066 280432 144154
rect 280540 144066 280720 144154
rect 280828 144066 281008 144154
rect 281116 144066 281296 144154
rect 281404 144066 281584 144154
rect 281692 144066 281872 144154
rect 281980 144066 282160 144154
rect 282414 144066 282594 144154
rect 282702 144066 282882 144154
rect 282990 144066 283170 144154
rect 283278 144066 283458 144154
rect 283566 144066 283746 144154
rect 283854 144066 284034 144154
rect 284142 144066 284322 144154
rect 284430 144066 284610 144154
rect 284864 144066 285044 144154
rect 285152 144066 285332 144154
rect 285440 144066 285620 144154
rect 285728 144066 285908 144154
rect 286016 144066 286196 144154
rect 286304 144066 286484 144154
rect 286592 144066 286772 144154
rect 286880 144066 287060 144154
rect 287314 144066 287494 144154
rect 287602 144066 287782 144154
rect 287890 144066 288070 144154
rect 288178 144066 288358 144154
rect 288466 144066 288646 144154
rect 288754 144066 288934 144154
rect 289042 144066 289222 144154
rect 289330 144066 289510 144154
rect 289764 144066 289944 144154
rect 290052 144066 290232 144154
rect 290340 144066 290520 144154
rect 290628 144066 290808 144154
rect 290916 144066 291096 144154
rect 291204 144066 291384 144154
rect 291492 144066 291672 144154
rect 291780 144066 291960 144154
rect 292214 144066 292394 144154
rect 292502 144066 292682 144154
rect 292790 144066 292970 144154
rect 293078 144066 293258 144154
rect 293366 144066 293546 144154
rect 293654 144066 293834 144154
rect 293942 144066 294122 144154
rect 294230 144066 294410 144154
rect 294664 144066 294844 144154
rect 294952 144066 295132 144154
rect 295240 144066 295420 144154
rect 295528 144066 295708 144154
rect 295816 144066 295996 144154
rect 296104 144066 296284 144154
rect 296392 144066 296572 144154
rect 296680 144066 296860 144154
rect 297114 144066 297294 144154
rect 297402 144066 297582 144154
rect 297690 144066 297870 144154
rect 297978 144066 298158 144154
rect 298266 144066 298446 144154
rect 298554 144066 298734 144154
rect 298842 144066 299022 144154
rect 299130 144066 299310 144154
rect 299564 144066 299744 144154
rect 299852 144066 300032 144154
rect 300140 144066 300320 144154
rect 300428 144066 300608 144154
rect 300716 144066 300896 144154
rect 301004 144066 301184 144154
rect 301292 144066 301472 144154
rect 301580 144066 301760 144154
rect 302014 144066 302194 144154
rect 302302 144066 302482 144154
rect 302590 144066 302770 144154
rect 302878 144066 303058 144154
rect 303166 144066 303346 144154
rect 303454 144066 303634 144154
rect 303742 144066 303922 144154
rect 304030 144066 304210 144154
rect 304464 144066 304644 144154
rect 304752 144066 304932 144154
rect 305040 144066 305220 144154
rect 305328 144066 305508 144154
rect 305616 144066 305796 144154
rect 305904 144066 306084 144154
rect 306192 144066 306372 144154
rect 306480 144066 306660 144154
rect 306914 144066 307094 144154
rect 307202 144066 307382 144154
rect 307490 144066 307670 144154
rect 307778 144066 307958 144154
rect 308066 144066 308246 144154
rect 308354 144066 308534 144154
rect 308642 144066 308822 144154
rect 308930 144066 309110 144154
rect 309364 144066 309544 144154
rect 309652 144066 309832 144154
rect 309940 144066 310120 144154
rect 310228 144066 310408 144154
rect 310516 144066 310696 144154
rect 310804 144066 310984 144154
rect 311092 144066 311272 144154
rect 311380 144066 311560 144154
rect 311814 144066 311994 144154
rect 312102 144066 312282 144154
rect 312390 144066 312570 144154
rect 312678 144066 312858 144154
rect 312966 144066 313146 144154
rect 313254 144066 313434 144154
rect 313542 144066 313722 144154
rect 313830 144066 314010 144154
rect 314264 144066 314444 144154
rect 314552 144066 314732 144154
rect 314840 144066 315020 144154
rect 315128 144066 315308 144154
rect 315416 144066 315596 144154
rect 315704 144066 315884 144154
rect 315992 144066 316172 144154
rect 316280 144066 316460 144154
rect 316714 144066 316894 144154
rect 317002 144066 317182 144154
rect 317290 144066 317470 144154
rect 317578 144066 317758 144154
rect 317866 144066 318046 144154
rect 318154 144066 318334 144154
rect 318442 144066 318622 144154
rect 318730 144066 318910 144154
rect 319164 144066 319344 144154
rect 319452 144066 319632 144154
rect 319740 144066 319920 144154
rect 320028 144066 320208 144154
rect 320316 144066 320496 144154
rect 320604 144066 320784 144154
rect 320892 144066 321072 144154
rect 321180 144066 321360 144154
rect 321614 144066 321794 144154
rect 321902 144066 322082 144154
rect 322190 144066 322370 144154
rect 322478 144066 322658 144154
rect 322766 144066 322946 144154
rect 323054 144066 323234 144154
rect 323342 144066 323522 144154
rect 323630 144066 323810 144154
rect 324064 144066 324244 144154
rect 324352 144066 324532 144154
rect 324640 144066 324820 144154
rect 324928 144066 325108 144154
rect 325216 144066 325396 144154
rect 325504 144066 325684 144154
rect 325792 144066 325972 144154
rect 326080 144066 326260 144154
rect 326514 144066 326694 144154
rect 326802 144066 326982 144154
rect 327090 144066 327270 144154
rect 327378 144066 327558 144154
rect 327666 144066 327846 144154
rect 327954 144066 328134 144154
rect 328242 144066 328422 144154
rect 328530 144066 328710 144154
rect 328964 144066 329144 144154
rect 329252 144066 329432 144154
rect 329540 144066 329720 144154
rect 329828 144066 330008 144154
rect 330116 144066 330296 144154
rect 330404 144066 330584 144154
rect 330692 144066 330872 144154
rect 330980 144066 331160 144154
rect 331414 144066 331594 144154
rect 331702 144066 331882 144154
rect 331990 144066 332170 144154
rect 332278 144066 332458 144154
rect 332566 144066 332746 144154
rect 332854 144066 333034 144154
rect 333142 144066 333322 144154
rect 333430 144066 333610 144154
rect 333864 144066 334044 144154
rect 334152 144066 334332 144154
rect 334440 144066 334620 144154
rect 334728 144066 334908 144154
rect 335016 144066 335196 144154
rect 335304 144066 335484 144154
rect 335592 144066 335772 144154
rect 335880 144066 336060 144154
rect 336314 144066 336494 144154
rect 336602 144066 336782 144154
rect 336890 144066 337070 144154
rect 337178 144066 337358 144154
rect 337466 144066 337646 144154
rect 337754 144066 337934 144154
rect 338042 144066 338222 144154
rect 338330 144066 338510 144154
rect 338764 144066 338944 144154
rect 339052 144066 339232 144154
rect 339340 144066 339520 144154
rect 339628 144066 339808 144154
rect 339916 144066 340096 144154
rect 340204 144066 340384 144154
rect 340492 144066 340672 144154
rect 340780 144066 340960 144154
rect 341214 144066 341394 144154
rect 341502 144066 341682 144154
rect 341790 144066 341970 144154
rect 342078 144066 342258 144154
rect 342366 144066 342546 144154
rect 342654 144066 342834 144154
rect 342942 144066 343122 144154
rect 343230 144066 343410 144154
rect 343664 144066 343844 144154
rect 343952 144066 344132 144154
rect 344240 144066 344420 144154
rect 344528 144066 344708 144154
rect 344816 144066 344996 144154
rect 345104 144066 345284 144154
rect 345392 144066 345572 144154
rect 345680 144066 345860 144154
rect 346114 144066 346294 144154
rect 346402 144066 346582 144154
rect 346690 144066 346870 144154
rect 346978 144066 347158 144154
rect 347266 144066 347446 144154
rect 347554 144066 347734 144154
rect 347842 144066 348022 144154
rect 348130 144066 348310 144154
rect 348564 144066 348744 144154
rect 348852 144066 349032 144154
rect 349140 144066 349320 144154
rect 349428 144066 349608 144154
rect 349716 144066 349896 144154
rect 350004 144066 350184 144154
rect 350292 144066 350472 144154
rect 350580 144066 350760 144154
rect 351014 144066 351194 144154
rect 351302 144066 351482 144154
rect 351590 144066 351770 144154
rect 351878 144066 352058 144154
rect 352166 144066 352346 144154
rect 352454 144066 352634 144154
rect 352742 144066 352922 144154
rect 353030 144066 353210 144154
rect 353464 144066 353644 144154
rect 353752 144066 353932 144154
rect 354040 144066 354220 144154
rect 354328 144066 354508 144154
rect 354616 144066 354796 144154
rect 354904 144066 355084 144154
rect 355192 144066 355372 144154
rect 355480 144066 355660 144154
rect 355914 144066 356094 144154
rect 356202 144066 356382 144154
rect 356490 144066 356670 144154
rect 356778 144066 356958 144154
rect 357066 144066 357246 144154
rect 357354 144066 357534 144154
rect 357642 144066 357822 144154
rect 357930 144066 358110 144154
rect 358364 144066 358544 144154
rect 358652 144066 358832 144154
rect 358940 144066 359120 144154
rect 359228 144066 359408 144154
rect 359516 144066 359696 144154
rect 359804 144066 359984 144154
rect 360092 144066 360272 144154
rect 360380 144066 360560 144154
rect 360814 144066 360994 144154
rect 361102 144066 361282 144154
rect 361390 144066 361570 144154
rect 361678 144066 361858 144154
rect 361966 144066 362146 144154
rect 362254 144066 362434 144154
rect 362542 144066 362722 144154
rect 362830 144066 363010 144154
rect 363264 144066 363444 144154
rect 363552 144066 363732 144154
rect 363840 144066 364020 144154
rect 364128 144066 364308 144154
rect 364416 144066 364596 144154
rect 364704 144066 364884 144154
rect 364992 144066 365172 144154
rect 365280 144066 365460 144154
rect 365714 144066 365894 144154
rect 366002 144066 366182 144154
rect 366290 144066 366470 144154
rect 366578 144066 366758 144154
rect 366866 144066 367046 144154
rect 367154 144066 367334 144154
rect 367442 144066 367622 144154
rect 367730 144066 367910 144154
rect 243214 143590 243394 143678
rect 243502 143590 243682 143678
rect 243790 143590 243970 143678
rect 244078 143590 244258 143678
rect 244366 143590 244546 143678
rect 244654 143590 244834 143678
rect 244942 143590 245122 143678
rect 245230 143590 245410 143678
rect 245664 143590 245844 143678
rect 245952 143590 246132 143678
rect 246240 143590 246420 143678
rect 246528 143590 246708 143678
rect 246816 143590 246996 143678
rect 247104 143590 247284 143678
rect 247392 143590 247572 143678
rect 247680 143590 247860 143678
rect 248114 143590 248294 143678
rect 248402 143590 248582 143678
rect 248690 143590 248870 143678
rect 248978 143590 249158 143678
rect 249266 143590 249446 143678
rect 249554 143590 249734 143678
rect 249842 143590 250022 143678
rect 250130 143590 250310 143678
rect 250564 143590 250744 143678
rect 250852 143590 251032 143678
rect 251140 143590 251320 143678
rect 251428 143590 251608 143678
rect 251716 143590 251896 143678
rect 252004 143590 252184 143678
rect 252292 143590 252472 143678
rect 252580 143590 252760 143678
rect 253014 143590 253194 143678
rect 253302 143590 253482 143678
rect 253590 143590 253770 143678
rect 253878 143590 254058 143678
rect 254166 143590 254346 143678
rect 254454 143590 254634 143678
rect 254742 143590 254922 143678
rect 255030 143590 255210 143678
rect 255464 143590 255644 143678
rect 255752 143590 255932 143678
rect 256040 143590 256220 143678
rect 256328 143590 256508 143678
rect 256616 143590 256796 143678
rect 256904 143590 257084 143678
rect 257192 143590 257372 143678
rect 257480 143590 257660 143678
rect 257914 143590 258094 143678
rect 258202 143590 258382 143678
rect 258490 143590 258670 143678
rect 258778 143590 258958 143678
rect 259066 143590 259246 143678
rect 259354 143590 259534 143678
rect 259642 143590 259822 143678
rect 259930 143590 260110 143678
rect 260364 143590 260544 143678
rect 260652 143590 260832 143678
rect 260940 143590 261120 143678
rect 261228 143590 261408 143678
rect 261516 143590 261696 143678
rect 261804 143590 261984 143678
rect 262092 143590 262272 143678
rect 262380 143590 262560 143678
rect 262814 143590 262994 143678
rect 263102 143590 263282 143678
rect 263390 143590 263570 143678
rect 263678 143590 263858 143678
rect 263966 143590 264146 143678
rect 264254 143590 264434 143678
rect 264542 143590 264722 143678
rect 264830 143590 265010 143678
rect 265264 143590 265444 143678
rect 265552 143590 265732 143678
rect 265840 143590 266020 143678
rect 266128 143590 266308 143678
rect 266416 143590 266596 143678
rect 266704 143590 266884 143678
rect 266992 143590 267172 143678
rect 267280 143590 267460 143678
rect 267714 143590 267894 143678
rect 268002 143590 268182 143678
rect 268290 143590 268470 143678
rect 268578 143590 268758 143678
rect 268866 143590 269046 143678
rect 269154 143590 269334 143678
rect 269442 143590 269622 143678
rect 269730 143590 269910 143678
rect 270164 143590 270344 143678
rect 270452 143590 270632 143678
rect 270740 143590 270920 143678
rect 271028 143590 271208 143678
rect 271316 143590 271496 143678
rect 271604 143590 271784 143678
rect 271892 143590 272072 143678
rect 272180 143590 272360 143678
rect 272614 143590 272794 143678
rect 272902 143590 273082 143678
rect 273190 143590 273370 143678
rect 273478 143590 273658 143678
rect 273766 143590 273946 143678
rect 274054 143590 274234 143678
rect 274342 143590 274522 143678
rect 274630 143590 274810 143678
rect 275064 143590 275244 143678
rect 275352 143590 275532 143678
rect 275640 143590 275820 143678
rect 275928 143590 276108 143678
rect 276216 143590 276396 143678
rect 276504 143590 276684 143678
rect 276792 143590 276972 143678
rect 277080 143590 277260 143678
rect 277514 143590 277694 143678
rect 277802 143590 277982 143678
rect 278090 143590 278270 143678
rect 278378 143590 278558 143678
rect 278666 143590 278846 143678
rect 278954 143590 279134 143678
rect 279242 143590 279422 143678
rect 279530 143590 279710 143678
rect 279964 143590 280144 143678
rect 280252 143590 280432 143678
rect 280540 143590 280720 143678
rect 280828 143590 281008 143678
rect 281116 143590 281296 143678
rect 281404 143590 281584 143678
rect 281692 143590 281872 143678
rect 281980 143590 282160 143678
rect 282414 143590 282594 143678
rect 282702 143590 282882 143678
rect 282990 143590 283170 143678
rect 283278 143590 283458 143678
rect 283566 143590 283746 143678
rect 283854 143590 284034 143678
rect 284142 143590 284322 143678
rect 284430 143590 284610 143678
rect 284864 143590 285044 143678
rect 285152 143590 285332 143678
rect 285440 143590 285620 143678
rect 285728 143590 285908 143678
rect 286016 143590 286196 143678
rect 286304 143590 286484 143678
rect 286592 143590 286772 143678
rect 286880 143590 287060 143678
rect 287314 143590 287494 143678
rect 287602 143590 287782 143678
rect 287890 143590 288070 143678
rect 288178 143590 288358 143678
rect 288466 143590 288646 143678
rect 288754 143590 288934 143678
rect 289042 143590 289222 143678
rect 289330 143590 289510 143678
rect 289764 143590 289944 143678
rect 290052 143590 290232 143678
rect 290340 143590 290520 143678
rect 290628 143590 290808 143678
rect 290916 143590 291096 143678
rect 291204 143590 291384 143678
rect 291492 143590 291672 143678
rect 291780 143590 291960 143678
rect 292214 143590 292394 143678
rect 292502 143590 292682 143678
rect 292790 143590 292970 143678
rect 293078 143590 293258 143678
rect 293366 143590 293546 143678
rect 293654 143590 293834 143678
rect 293942 143590 294122 143678
rect 294230 143590 294410 143678
rect 294664 143590 294844 143678
rect 294952 143590 295132 143678
rect 295240 143590 295420 143678
rect 295528 143590 295708 143678
rect 295816 143590 295996 143678
rect 296104 143590 296284 143678
rect 296392 143590 296572 143678
rect 296680 143590 296860 143678
rect 297114 143590 297294 143678
rect 297402 143590 297582 143678
rect 297690 143590 297870 143678
rect 297978 143590 298158 143678
rect 298266 143590 298446 143678
rect 298554 143590 298734 143678
rect 298842 143590 299022 143678
rect 299130 143590 299310 143678
rect 299564 143590 299744 143678
rect 299852 143590 300032 143678
rect 300140 143590 300320 143678
rect 300428 143590 300608 143678
rect 300716 143590 300896 143678
rect 301004 143590 301184 143678
rect 301292 143590 301472 143678
rect 301580 143590 301760 143678
rect 302014 143590 302194 143678
rect 302302 143590 302482 143678
rect 302590 143590 302770 143678
rect 302878 143590 303058 143678
rect 303166 143590 303346 143678
rect 303454 143590 303634 143678
rect 303742 143590 303922 143678
rect 304030 143590 304210 143678
rect 304464 143590 304644 143678
rect 304752 143590 304932 143678
rect 305040 143590 305220 143678
rect 305328 143590 305508 143678
rect 305616 143590 305796 143678
rect 305904 143590 306084 143678
rect 306192 143590 306372 143678
rect 306480 143590 306660 143678
rect 306914 143590 307094 143678
rect 307202 143590 307382 143678
rect 307490 143590 307670 143678
rect 307778 143590 307958 143678
rect 308066 143590 308246 143678
rect 308354 143590 308534 143678
rect 308642 143590 308822 143678
rect 308930 143590 309110 143678
rect 309364 143590 309544 143678
rect 309652 143590 309832 143678
rect 309940 143590 310120 143678
rect 310228 143590 310408 143678
rect 310516 143590 310696 143678
rect 310804 143590 310984 143678
rect 311092 143590 311272 143678
rect 311380 143590 311560 143678
rect 311814 143590 311994 143678
rect 312102 143590 312282 143678
rect 312390 143590 312570 143678
rect 312678 143590 312858 143678
rect 312966 143590 313146 143678
rect 313254 143590 313434 143678
rect 313542 143590 313722 143678
rect 313830 143590 314010 143678
rect 314264 143590 314444 143678
rect 314552 143590 314732 143678
rect 314840 143590 315020 143678
rect 315128 143590 315308 143678
rect 315416 143590 315596 143678
rect 315704 143590 315884 143678
rect 315992 143590 316172 143678
rect 316280 143590 316460 143678
rect 316714 143590 316894 143678
rect 317002 143590 317182 143678
rect 317290 143590 317470 143678
rect 317578 143590 317758 143678
rect 317866 143590 318046 143678
rect 318154 143590 318334 143678
rect 318442 143590 318622 143678
rect 318730 143590 318910 143678
rect 319164 143590 319344 143678
rect 319452 143590 319632 143678
rect 319740 143590 319920 143678
rect 320028 143590 320208 143678
rect 320316 143590 320496 143678
rect 320604 143590 320784 143678
rect 320892 143590 321072 143678
rect 321180 143590 321360 143678
rect 321614 143590 321794 143678
rect 321902 143590 322082 143678
rect 322190 143590 322370 143678
rect 322478 143590 322658 143678
rect 322766 143590 322946 143678
rect 323054 143590 323234 143678
rect 323342 143590 323522 143678
rect 323630 143590 323810 143678
rect 324064 143590 324244 143678
rect 324352 143590 324532 143678
rect 324640 143590 324820 143678
rect 324928 143590 325108 143678
rect 325216 143590 325396 143678
rect 325504 143590 325684 143678
rect 325792 143590 325972 143678
rect 326080 143590 326260 143678
rect 326514 143590 326694 143678
rect 326802 143590 326982 143678
rect 327090 143590 327270 143678
rect 327378 143590 327558 143678
rect 327666 143590 327846 143678
rect 327954 143590 328134 143678
rect 328242 143590 328422 143678
rect 328530 143590 328710 143678
rect 328964 143590 329144 143678
rect 329252 143590 329432 143678
rect 329540 143590 329720 143678
rect 329828 143590 330008 143678
rect 330116 143590 330296 143678
rect 330404 143590 330584 143678
rect 330692 143590 330872 143678
rect 330980 143590 331160 143678
rect 331414 143590 331594 143678
rect 331702 143590 331882 143678
rect 331990 143590 332170 143678
rect 332278 143590 332458 143678
rect 332566 143590 332746 143678
rect 332854 143590 333034 143678
rect 333142 143590 333322 143678
rect 333430 143590 333610 143678
rect 333864 143590 334044 143678
rect 334152 143590 334332 143678
rect 334440 143590 334620 143678
rect 334728 143590 334908 143678
rect 335016 143590 335196 143678
rect 335304 143590 335484 143678
rect 335592 143590 335772 143678
rect 335880 143590 336060 143678
rect 336314 143590 336494 143678
rect 336602 143590 336782 143678
rect 336890 143590 337070 143678
rect 337178 143590 337358 143678
rect 337466 143590 337646 143678
rect 337754 143590 337934 143678
rect 338042 143590 338222 143678
rect 338330 143590 338510 143678
rect 338764 143590 338944 143678
rect 339052 143590 339232 143678
rect 339340 143590 339520 143678
rect 339628 143590 339808 143678
rect 339916 143590 340096 143678
rect 340204 143590 340384 143678
rect 340492 143590 340672 143678
rect 340780 143590 340960 143678
rect 341214 143590 341394 143678
rect 341502 143590 341682 143678
rect 341790 143590 341970 143678
rect 342078 143590 342258 143678
rect 342366 143590 342546 143678
rect 342654 143590 342834 143678
rect 342942 143590 343122 143678
rect 343230 143590 343410 143678
rect 343664 143590 343844 143678
rect 343952 143590 344132 143678
rect 344240 143590 344420 143678
rect 344528 143590 344708 143678
rect 344816 143590 344996 143678
rect 345104 143590 345284 143678
rect 345392 143590 345572 143678
rect 345680 143590 345860 143678
rect 346114 143590 346294 143678
rect 346402 143590 346582 143678
rect 346690 143590 346870 143678
rect 346978 143590 347158 143678
rect 347266 143590 347446 143678
rect 347554 143590 347734 143678
rect 347842 143590 348022 143678
rect 348130 143590 348310 143678
rect 348564 143590 348744 143678
rect 348852 143590 349032 143678
rect 349140 143590 349320 143678
rect 349428 143590 349608 143678
rect 349716 143590 349896 143678
rect 350004 143590 350184 143678
rect 350292 143590 350472 143678
rect 350580 143590 350760 143678
rect 351014 143590 351194 143678
rect 351302 143590 351482 143678
rect 351590 143590 351770 143678
rect 351878 143590 352058 143678
rect 352166 143590 352346 143678
rect 352454 143590 352634 143678
rect 352742 143590 352922 143678
rect 353030 143590 353210 143678
rect 353464 143590 353644 143678
rect 353752 143590 353932 143678
rect 354040 143590 354220 143678
rect 354328 143590 354508 143678
rect 354616 143590 354796 143678
rect 354904 143590 355084 143678
rect 355192 143590 355372 143678
rect 355480 143590 355660 143678
rect 355914 143590 356094 143678
rect 356202 143590 356382 143678
rect 356490 143590 356670 143678
rect 356778 143590 356958 143678
rect 357066 143590 357246 143678
rect 357354 143590 357534 143678
rect 357642 143590 357822 143678
rect 357930 143590 358110 143678
rect 358364 143590 358544 143678
rect 358652 143590 358832 143678
rect 358940 143590 359120 143678
rect 359228 143590 359408 143678
rect 359516 143590 359696 143678
rect 359804 143590 359984 143678
rect 360092 143590 360272 143678
rect 360380 143590 360560 143678
rect 360814 143590 360994 143678
rect 361102 143590 361282 143678
rect 361390 143590 361570 143678
rect 361678 143590 361858 143678
rect 361966 143590 362146 143678
rect 362254 143590 362434 143678
rect 362542 143590 362722 143678
rect 362830 143590 363010 143678
rect 363264 143590 363444 143678
rect 363552 143590 363732 143678
rect 363840 143590 364020 143678
rect 364128 143590 364308 143678
rect 364416 143590 364596 143678
rect 364704 143590 364884 143678
rect 364992 143590 365172 143678
rect 365280 143590 365460 143678
rect 365714 143590 365894 143678
rect 366002 143590 366182 143678
rect 366290 143590 366470 143678
rect 366578 143590 366758 143678
rect 366866 143590 367046 143678
rect 367154 143590 367334 143678
rect 367442 143590 367622 143678
rect 367730 143590 367910 143678
rect 243214 143374 243394 143462
rect 243502 143374 243682 143462
rect 243790 143374 243970 143462
rect 244078 143374 244258 143462
rect 244366 143374 244546 143462
rect 244654 143374 244834 143462
rect 244942 143374 245122 143462
rect 245230 143374 245410 143462
rect 245664 143374 245844 143462
rect 245952 143374 246132 143462
rect 246240 143374 246420 143462
rect 246528 143374 246708 143462
rect 246816 143374 246996 143462
rect 247104 143374 247284 143462
rect 247392 143374 247572 143462
rect 247680 143374 247860 143462
rect 248114 143374 248294 143462
rect 248402 143374 248582 143462
rect 248690 143374 248870 143462
rect 248978 143374 249158 143462
rect 249266 143374 249446 143462
rect 249554 143374 249734 143462
rect 249842 143374 250022 143462
rect 250130 143374 250310 143462
rect 250564 143374 250744 143462
rect 250852 143374 251032 143462
rect 251140 143374 251320 143462
rect 251428 143374 251608 143462
rect 251716 143374 251896 143462
rect 252004 143374 252184 143462
rect 252292 143374 252472 143462
rect 252580 143374 252760 143462
rect 253014 143374 253194 143462
rect 253302 143374 253482 143462
rect 253590 143374 253770 143462
rect 253878 143374 254058 143462
rect 254166 143374 254346 143462
rect 254454 143374 254634 143462
rect 254742 143374 254922 143462
rect 255030 143374 255210 143462
rect 255464 143374 255644 143462
rect 255752 143374 255932 143462
rect 256040 143374 256220 143462
rect 256328 143374 256508 143462
rect 256616 143374 256796 143462
rect 256904 143374 257084 143462
rect 257192 143374 257372 143462
rect 257480 143374 257660 143462
rect 257914 143374 258094 143462
rect 258202 143374 258382 143462
rect 258490 143374 258670 143462
rect 258778 143374 258958 143462
rect 259066 143374 259246 143462
rect 259354 143374 259534 143462
rect 259642 143374 259822 143462
rect 259930 143374 260110 143462
rect 260364 143374 260544 143462
rect 260652 143374 260832 143462
rect 260940 143374 261120 143462
rect 261228 143374 261408 143462
rect 261516 143374 261696 143462
rect 261804 143374 261984 143462
rect 262092 143374 262272 143462
rect 262380 143374 262560 143462
rect 262814 143374 262994 143462
rect 263102 143374 263282 143462
rect 263390 143374 263570 143462
rect 263678 143374 263858 143462
rect 263966 143374 264146 143462
rect 264254 143374 264434 143462
rect 264542 143374 264722 143462
rect 264830 143374 265010 143462
rect 265264 143374 265444 143462
rect 265552 143374 265732 143462
rect 265840 143374 266020 143462
rect 266128 143374 266308 143462
rect 266416 143374 266596 143462
rect 266704 143374 266884 143462
rect 266992 143374 267172 143462
rect 267280 143374 267460 143462
rect 267714 143374 267894 143462
rect 268002 143374 268182 143462
rect 268290 143374 268470 143462
rect 268578 143374 268758 143462
rect 268866 143374 269046 143462
rect 269154 143374 269334 143462
rect 269442 143374 269622 143462
rect 269730 143374 269910 143462
rect 270164 143374 270344 143462
rect 270452 143374 270632 143462
rect 270740 143374 270920 143462
rect 271028 143374 271208 143462
rect 271316 143374 271496 143462
rect 271604 143374 271784 143462
rect 271892 143374 272072 143462
rect 272180 143374 272360 143462
rect 272614 143374 272794 143462
rect 272902 143374 273082 143462
rect 273190 143374 273370 143462
rect 273478 143374 273658 143462
rect 273766 143374 273946 143462
rect 274054 143374 274234 143462
rect 274342 143374 274522 143462
rect 274630 143374 274810 143462
rect 275064 143374 275244 143462
rect 275352 143374 275532 143462
rect 275640 143374 275820 143462
rect 275928 143374 276108 143462
rect 276216 143374 276396 143462
rect 276504 143374 276684 143462
rect 276792 143374 276972 143462
rect 277080 143374 277260 143462
rect 277514 143374 277694 143462
rect 277802 143374 277982 143462
rect 278090 143374 278270 143462
rect 278378 143374 278558 143462
rect 278666 143374 278846 143462
rect 278954 143374 279134 143462
rect 279242 143374 279422 143462
rect 279530 143374 279710 143462
rect 279964 143374 280144 143462
rect 280252 143374 280432 143462
rect 280540 143374 280720 143462
rect 280828 143374 281008 143462
rect 281116 143374 281296 143462
rect 281404 143374 281584 143462
rect 281692 143374 281872 143462
rect 281980 143374 282160 143462
rect 282414 143374 282594 143462
rect 282702 143374 282882 143462
rect 282990 143374 283170 143462
rect 283278 143374 283458 143462
rect 283566 143374 283746 143462
rect 283854 143374 284034 143462
rect 284142 143374 284322 143462
rect 284430 143374 284610 143462
rect 284864 143374 285044 143462
rect 285152 143374 285332 143462
rect 285440 143374 285620 143462
rect 285728 143374 285908 143462
rect 286016 143374 286196 143462
rect 286304 143374 286484 143462
rect 286592 143374 286772 143462
rect 286880 143374 287060 143462
rect 287314 143374 287494 143462
rect 287602 143374 287782 143462
rect 287890 143374 288070 143462
rect 288178 143374 288358 143462
rect 288466 143374 288646 143462
rect 288754 143374 288934 143462
rect 289042 143374 289222 143462
rect 289330 143374 289510 143462
rect 289764 143374 289944 143462
rect 290052 143374 290232 143462
rect 290340 143374 290520 143462
rect 290628 143374 290808 143462
rect 290916 143374 291096 143462
rect 291204 143374 291384 143462
rect 291492 143374 291672 143462
rect 291780 143374 291960 143462
rect 292214 143374 292394 143462
rect 292502 143374 292682 143462
rect 292790 143374 292970 143462
rect 293078 143374 293258 143462
rect 293366 143374 293546 143462
rect 293654 143374 293834 143462
rect 293942 143374 294122 143462
rect 294230 143374 294410 143462
rect 294664 143374 294844 143462
rect 294952 143374 295132 143462
rect 295240 143374 295420 143462
rect 295528 143374 295708 143462
rect 295816 143374 295996 143462
rect 296104 143374 296284 143462
rect 296392 143374 296572 143462
rect 296680 143374 296860 143462
rect 297114 143374 297294 143462
rect 297402 143374 297582 143462
rect 297690 143374 297870 143462
rect 297978 143374 298158 143462
rect 298266 143374 298446 143462
rect 298554 143374 298734 143462
rect 298842 143374 299022 143462
rect 299130 143374 299310 143462
rect 299564 143374 299744 143462
rect 299852 143374 300032 143462
rect 300140 143374 300320 143462
rect 300428 143374 300608 143462
rect 300716 143374 300896 143462
rect 301004 143374 301184 143462
rect 301292 143374 301472 143462
rect 301580 143374 301760 143462
rect 302014 143374 302194 143462
rect 302302 143374 302482 143462
rect 302590 143374 302770 143462
rect 302878 143374 303058 143462
rect 303166 143374 303346 143462
rect 303454 143374 303634 143462
rect 303742 143374 303922 143462
rect 304030 143374 304210 143462
rect 304464 143374 304644 143462
rect 304752 143374 304932 143462
rect 305040 143374 305220 143462
rect 305328 143374 305508 143462
rect 305616 143374 305796 143462
rect 305904 143374 306084 143462
rect 306192 143374 306372 143462
rect 306480 143374 306660 143462
rect 306914 143374 307094 143462
rect 307202 143374 307382 143462
rect 307490 143374 307670 143462
rect 307778 143374 307958 143462
rect 308066 143374 308246 143462
rect 308354 143374 308534 143462
rect 308642 143374 308822 143462
rect 308930 143374 309110 143462
rect 309364 143374 309544 143462
rect 309652 143374 309832 143462
rect 309940 143374 310120 143462
rect 310228 143374 310408 143462
rect 310516 143374 310696 143462
rect 310804 143374 310984 143462
rect 311092 143374 311272 143462
rect 311380 143374 311560 143462
rect 311814 143374 311994 143462
rect 312102 143374 312282 143462
rect 312390 143374 312570 143462
rect 312678 143374 312858 143462
rect 312966 143374 313146 143462
rect 313254 143374 313434 143462
rect 313542 143374 313722 143462
rect 313830 143374 314010 143462
rect 314264 143374 314444 143462
rect 314552 143374 314732 143462
rect 314840 143374 315020 143462
rect 315128 143374 315308 143462
rect 315416 143374 315596 143462
rect 315704 143374 315884 143462
rect 315992 143374 316172 143462
rect 316280 143374 316460 143462
rect 316714 143374 316894 143462
rect 317002 143374 317182 143462
rect 317290 143374 317470 143462
rect 317578 143374 317758 143462
rect 317866 143374 318046 143462
rect 318154 143374 318334 143462
rect 318442 143374 318622 143462
rect 318730 143374 318910 143462
rect 319164 143374 319344 143462
rect 319452 143374 319632 143462
rect 319740 143374 319920 143462
rect 320028 143374 320208 143462
rect 320316 143374 320496 143462
rect 320604 143374 320784 143462
rect 320892 143374 321072 143462
rect 321180 143374 321360 143462
rect 321614 143374 321794 143462
rect 321902 143374 322082 143462
rect 322190 143374 322370 143462
rect 322478 143374 322658 143462
rect 322766 143374 322946 143462
rect 323054 143374 323234 143462
rect 323342 143374 323522 143462
rect 323630 143374 323810 143462
rect 324064 143374 324244 143462
rect 324352 143374 324532 143462
rect 324640 143374 324820 143462
rect 324928 143374 325108 143462
rect 325216 143374 325396 143462
rect 325504 143374 325684 143462
rect 325792 143374 325972 143462
rect 326080 143374 326260 143462
rect 326514 143374 326694 143462
rect 326802 143374 326982 143462
rect 327090 143374 327270 143462
rect 327378 143374 327558 143462
rect 327666 143374 327846 143462
rect 327954 143374 328134 143462
rect 328242 143374 328422 143462
rect 328530 143374 328710 143462
rect 328964 143374 329144 143462
rect 329252 143374 329432 143462
rect 329540 143374 329720 143462
rect 329828 143374 330008 143462
rect 330116 143374 330296 143462
rect 330404 143374 330584 143462
rect 330692 143374 330872 143462
rect 330980 143374 331160 143462
rect 331414 143374 331594 143462
rect 331702 143374 331882 143462
rect 331990 143374 332170 143462
rect 332278 143374 332458 143462
rect 332566 143374 332746 143462
rect 332854 143374 333034 143462
rect 333142 143374 333322 143462
rect 333430 143374 333610 143462
rect 333864 143374 334044 143462
rect 334152 143374 334332 143462
rect 334440 143374 334620 143462
rect 334728 143374 334908 143462
rect 335016 143374 335196 143462
rect 335304 143374 335484 143462
rect 335592 143374 335772 143462
rect 335880 143374 336060 143462
rect 336314 143374 336494 143462
rect 336602 143374 336782 143462
rect 336890 143374 337070 143462
rect 337178 143374 337358 143462
rect 337466 143374 337646 143462
rect 337754 143374 337934 143462
rect 338042 143374 338222 143462
rect 338330 143374 338510 143462
rect 338764 143374 338944 143462
rect 339052 143374 339232 143462
rect 339340 143374 339520 143462
rect 339628 143374 339808 143462
rect 339916 143374 340096 143462
rect 340204 143374 340384 143462
rect 340492 143374 340672 143462
rect 340780 143374 340960 143462
rect 341214 143374 341394 143462
rect 341502 143374 341682 143462
rect 341790 143374 341970 143462
rect 342078 143374 342258 143462
rect 342366 143374 342546 143462
rect 342654 143374 342834 143462
rect 342942 143374 343122 143462
rect 343230 143374 343410 143462
rect 343664 143374 343844 143462
rect 343952 143374 344132 143462
rect 344240 143374 344420 143462
rect 344528 143374 344708 143462
rect 344816 143374 344996 143462
rect 345104 143374 345284 143462
rect 345392 143374 345572 143462
rect 345680 143374 345860 143462
rect 346114 143374 346294 143462
rect 346402 143374 346582 143462
rect 346690 143374 346870 143462
rect 346978 143374 347158 143462
rect 347266 143374 347446 143462
rect 347554 143374 347734 143462
rect 347842 143374 348022 143462
rect 348130 143374 348310 143462
rect 348564 143374 348744 143462
rect 348852 143374 349032 143462
rect 349140 143374 349320 143462
rect 349428 143374 349608 143462
rect 349716 143374 349896 143462
rect 350004 143374 350184 143462
rect 350292 143374 350472 143462
rect 350580 143374 350760 143462
rect 351014 143374 351194 143462
rect 351302 143374 351482 143462
rect 351590 143374 351770 143462
rect 351878 143374 352058 143462
rect 352166 143374 352346 143462
rect 352454 143374 352634 143462
rect 352742 143374 352922 143462
rect 353030 143374 353210 143462
rect 353464 143374 353644 143462
rect 353752 143374 353932 143462
rect 354040 143374 354220 143462
rect 354328 143374 354508 143462
rect 354616 143374 354796 143462
rect 354904 143374 355084 143462
rect 355192 143374 355372 143462
rect 355480 143374 355660 143462
rect 355914 143374 356094 143462
rect 356202 143374 356382 143462
rect 356490 143374 356670 143462
rect 356778 143374 356958 143462
rect 357066 143374 357246 143462
rect 357354 143374 357534 143462
rect 357642 143374 357822 143462
rect 357930 143374 358110 143462
rect 358364 143374 358544 143462
rect 358652 143374 358832 143462
rect 358940 143374 359120 143462
rect 359228 143374 359408 143462
rect 359516 143374 359696 143462
rect 359804 143374 359984 143462
rect 360092 143374 360272 143462
rect 360380 143374 360560 143462
rect 360814 143374 360994 143462
rect 361102 143374 361282 143462
rect 361390 143374 361570 143462
rect 361678 143374 361858 143462
rect 361966 143374 362146 143462
rect 362254 143374 362434 143462
rect 362542 143374 362722 143462
rect 362830 143374 363010 143462
rect 363264 143374 363444 143462
rect 363552 143374 363732 143462
rect 363840 143374 364020 143462
rect 364128 143374 364308 143462
rect 364416 143374 364596 143462
rect 364704 143374 364884 143462
rect 364992 143374 365172 143462
rect 365280 143374 365460 143462
rect 365714 143374 365894 143462
rect 366002 143374 366182 143462
rect 366290 143374 366470 143462
rect 366578 143374 366758 143462
rect 366866 143374 367046 143462
rect 367154 143374 367334 143462
rect 367442 143374 367622 143462
rect 367730 143374 367910 143462
rect 243214 142898 243394 142986
rect 243502 142898 243682 142986
rect 243790 142898 243970 142986
rect 244078 142898 244258 142986
rect 244366 142898 244546 142986
rect 244654 142898 244834 142986
rect 244942 142898 245122 142986
rect 245230 142898 245410 142986
rect 245664 142898 245844 142986
rect 245952 142898 246132 142986
rect 246240 142898 246420 142986
rect 246528 142898 246708 142986
rect 246816 142898 246996 142986
rect 247104 142898 247284 142986
rect 247392 142898 247572 142986
rect 247680 142898 247860 142986
rect 248114 142898 248294 142986
rect 248402 142898 248582 142986
rect 248690 142898 248870 142986
rect 248978 142898 249158 142986
rect 249266 142898 249446 142986
rect 249554 142898 249734 142986
rect 249842 142898 250022 142986
rect 250130 142898 250310 142986
rect 250564 142898 250744 142986
rect 250852 142898 251032 142986
rect 251140 142898 251320 142986
rect 251428 142898 251608 142986
rect 251716 142898 251896 142986
rect 252004 142898 252184 142986
rect 252292 142898 252472 142986
rect 252580 142898 252760 142986
rect 253014 142898 253194 142986
rect 253302 142898 253482 142986
rect 253590 142898 253770 142986
rect 253878 142898 254058 142986
rect 254166 142898 254346 142986
rect 254454 142898 254634 142986
rect 254742 142898 254922 142986
rect 255030 142898 255210 142986
rect 255464 142898 255644 142986
rect 255752 142898 255932 142986
rect 256040 142898 256220 142986
rect 256328 142898 256508 142986
rect 256616 142898 256796 142986
rect 256904 142898 257084 142986
rect 257192 142898 257372 142986
rect 257480 142898 257660 142986
rect 257914 142898 258094 142986
rect 258202 142898 258382 142986
rect 258490 142898 258670 142986
rect 258778 142898 258958 142986
rect 259066 142898 259246 142986
rect 259354 142898 259534 142986
rect 259642 142898 259822 142986
rect 259930 142898 260110 142986
rect 260364 142898 260544 142986
rect 260652 142898 260832 142986
rect 260940 142898 261120 142986
rect 261228 142898 261408 142986
rect 261516 142898 261696 142986
rect 261804 142898 261984 142986
rect 262092 142898 262272 142986
rect 262380 142898 262560 142986
rect 262814 142898 262994 142986
rect 263102 142898 263282 142986
rect 263390 142898 263570 142986
rect 263678 142898 263858 142986
rect 263966 142898 264146 142986
rect 264254 142898 264434 142986
rect 264542 142898 264722 142986
rect 264830 142898 265010 142986
rect 265264 142898 265444 142986
rect 265552 142898 265732 142986
rect 265840 142898 266020 142986
rect 266128 142898 266308 142986
rect 266416 142898 266596 142986
rect 266704 142898 266884 142986
rect 266992 142898 267172 142986
rect 267280 142898 267460 142986
rect 267714 142898 267894 142986
rect 268002 142898 268182 142986
rect 268290 142898 268470 142986
rect 268578 142898 268758 142986
rect 268866 142898 269046 142986
rect 269154 142898 269334 142986
rect 269442 142898 269622 142986
rect 269730 142898 269910 142986
rect 270164 142898 270344 142986
rect 270452 142898 270632 142986
rect 270740 142898 270920 142986
rect 271028 142898 271208 142986
rect 271316 142898 271496 142986
rect 271604 142898 271784 142986
rect 271892 142898 272072 142986
rect 272180 142898 272360 142986
rect 272614 142898 272794 142986
rect 272902 142898 273082 142986
rect 273190 142898 273370 142986
rect 273478 142898 273658 142986
rect 273766 142898 273946 142986
rect 274054 142898 274234 142986
rect 274342 142898 274522 142986
rect 274630 142898 274810 142986
rect 275064 142898 275244 142986
rect 275352 142898 275532 142986
rect 275640 142898 275820 142986
rect 275928 142898 276108 142986
rect 276216 142898 276396 142986
rect 276504 142898 276684 142986
rect 276792 142898 276972 142986
rect 277080 142898 277260 142986
rect 277514 142898 277694 142986
rect 277802 142898 277982 142986
rect 278090 142898 278270 142986
rect 278378 142898 278558 142986
rect 278666 142898 278846 142986
rect 278954 142898 279134 142986
rect 279242 142898 279422 142986
rect 279530 142898 279710 142986
rect 279964 142898 280144 142986
rect 280252 142898 280432 142986
rect 280540 142898 280720 142986
rect 280828 142898 281008 142986
rect 281116 142898 281296 142986
rect 281404 142898 281584 142986
rect 281692 142898 281872 142986
rect 281980 142898 282160 142986
rect 282414 142898 282594 142986
rect 282702 142898 282882 142986
rect 282990 142898 283170 142986
rect 283278 142898 283458 142986
rect 283566 142898 283746 142986
rect 283854 142898 284034 142986
rect 284142 142898 284322 142986
rect 284430 142898 284610 142986
rect 284864 142898 285044 142986
rect 285152 142898 285332 142986
rect 285440 142898 285620 142986
rect 285728 142898 285908 142986
rect 286016 142898 286196 142986
rect 286304 142898 286484 142986
rect 286592 142898 286772 142986
rect 286880 142898 287060 142986
rect 287314 142898 287494 142986
rect 287602 142898 287782 142986
rect 287890 142898 288070 142986
rect 288178 142898 288358 142986
rect 288466 142898 288646 142986
rect 288754 142898 288934 142986
rect 289042 142898 289222 142986
rect 289330 142898 289510 142986
rect 289764 142898 289944 142986
rect 290052 142898 290232 142986
rect 290340 142898 290520 142986
rect 290628 142898 290808 142986
rect 290916 142898 291096 142986
rect 291204 142898 291384 142986
rect 291492 142898 291672 142986
rect 291780 142898 291960 142986
rect 292214 142898 292394 142986
rect 292502 142898 292682 142986
rect 292790 142898 292970 142986
rect 293078 142898 293258 142986
rect 293366 142898 293546 142986
rect 293654 142898 293834 142986
rect 293942 142898 294122 142986
rect 294230 142898 294410 142986
rect 294664 142898 294844 142986
rect 294952 142898 295132 142986
rect 295240 142898 295420 142986
rect 295528 142898 295708 142986
rect 295816 142898 295996 142986
rect 296104 142898 296284 142986
rect 296392 142898 296572 142986
rect 296680 142898 296860 142986
rect 297114 142898 297294 142986
rect 297402 142898 297582 142986
rect 297690 142898 297870 142986
rect 297978 142898 298158 142986
rect 298266 142898 298446 142986
rect 298554 142898 298734 142986
rect 298842 142898 299022 142986
rect 299130 142898 299310 142986
rect 299564 142898 299744 142986
rect 299852 142898 300032 142986
rect 300140 142898 300320 142986
rect 300428 142898 300608 142986
rect 300716 142898 300896 142986
rect 301004 142898 301184 142986
rect 301292 142898 301472 142986
rect 301580 142898 301760 142986
rect 302014 142898 302194 142986
rect 302302 142898 302482 142986
rect 302590 142898 302770 142986
rect 302878 142898 303058 142986
rect 303166 142898 303346 142986
rect 303454 142898 303634 142986
rect 303742 142898 303922 142986
rect 304030 142898 304210 142986
rect 304464 142898 304644 142986
rect 304752 142898 304932 142986
rect 305040 142898 305220 142986
rect 305328 142898 305508 142986
rect 305616 142898 305796 142986
rect 305904 142898 306084 142986
rect 306192 142898 306372 142986
rect 306480 142898 306660 142986
rect 306914 142898 307094 142986
rect 307202 142898 307382 142986
rect 307490 142898 307670 142986
rect 307778 142898 307958 142986
rect 308066 142898 308246 142986
rect 308354 142898 308534 142986
rect 308642 142898 308822 142986
rect 308930 142898 309110 142986
rect 309364 142898 309544 142986
rect 309652 142898 309832 142986
rect 309940 142898 310120 142986
rect 310228 142898 310408 142986
rect 310516 142898 310696 142986
rect 310804 142898 310984 142986
rect 311092 142898 311272 142986
rect 311380 142898 311560 142986
rect 311814 142898 311994 142986
rect 312102 142898 312282 142986
rect 312390 142898 312570 142986
rect 312678 142898 312858 142986
rect 312966 142898 313146 142986
rect 313254 142898 313434 142986
rect 313542 142898 313722 142986
rect 313830 142898 314010 142986
rect 314264 142898 314444 142986
rect 314552 142898 314732 142986
rect 314840 142898 315020 142986
rect 315128 142898 315308 142986
rect 315416 142898 315596 142986
rect 315704 142898 315884 142986
rect 315992 142898 316172 142986
rect 316280 142898 316460 142986
rect 316714 142898 316894 142986
rect 317002 142898 317182 142986
rect 317290 142898 317470 142986
rect 317578 142898 317758 142986
rect 317866 142898 318046 142986
rect 318154 142898 318334 142986
rect 318442 142898 318622 142986
rect 318730 142898 318910 142986
rect 319164 142898 319344 142986
rect 319452 142898 319632 142986
rect 319740 142898 319920 142986
rect 320028 142898 320208 142986
rect 320316 142898 320496 142986
rect 320604 142898 320784 142986
rect 320892 142898 321072 142986
rect 321180 142898 321360 142986
rect 321614 142898 321794 142986
rect 321902 142898 322082 142986
rect 322190 142898 322370 142986
rect 322478 142898 322658 142986
rect 322766 142898 322946 142986
rect 323054 142898 323234 142986
rect 323342 142898 323522 142986
rect 323630 142898 323810 142986
rect 324064 142898 324244 142986
rect 324352 142898 324532 142986
rect 324640 142898 324820 142986
rect 324928 142898 325108 142986
rect 325216 142898 325396 142986
rect 325504 142898 325684 142986
rect 325792 142898 325972 142986
rect 326080 142898 326260 142986
rect 326514 142898 326694 142986
rect 326802 142898 326982 142986
rect 327090 142898 327270 142986
rect 327378 142898 327558 142986
rect 327666 142898 327846 142986
rect 327954 142898 328134 142986
rect 328242 142898 328422 142986
rect 328530 142898 328710 142986
rect 328964 142898 329144 142986
rect 329252 142898 329432 142986
rect 329540 142898 329720 142986
rect 329828 142898 330008 142986
rect 330116 142898 330296 142986
rect 330404 142898 330584 142986
rect 330692 142898 330872 142986
rect 330980 142898 331160 142986
rect 331414 142898 331594 142986
rect 331702 142898 331882 142986
rect 331990 142898 332170 142986
rect 332278 142898 332458 142986
rect 332566 142898 332746 142986
rect 332854 142898 333034 142986
rect 333142 142898 333322 142986
rect 333430 142898 333610 142986
rect 333864 142898 334044 142986
rect 334152 142898 334332 142986
rect 334440 142898 334620 142986
rect 334728 142898 334908 142986
rect 335016 142898 335196 142986
rect 335304 142898 335484 142986
rect 335592 142898 335772 142986
rect 335880 142898 336060 142986
rect 336314 142898 336494 142986
rect 336602 142898 336782 142986
rect 336890 142898 337070 142986
rect 337178 142898 337358 142986
rect 337466 142898 337646 142986
rect 337754 142898 337934 142986
rect 338042 142898 338222 142986
rect 338330 142898 338510 142986
rect 338764 142898 338944 142986
rect 339052 142898 339232 142986
rect 339340 142898 339520 142986
rect 339628 142898 339808 142986
rect 339916 142898 340096 142986
rect 340204 142898 340384 142986
rect 340492 142898 340672 142986
rect 340780 142898 340960 142986
rect 341214 142898 341394 142986
rect 341502 142898 341682 142986
rect 341790 142898 341970 142986
rect 342078 142898 342258 142986
rect 342366 142898 342546 142986
rect 342654 142898 342834 142986
rect 342942 142898 343122 142986
rect 343230 142898 343410 142986
rect 343664 142898 343844 142986
rect 343952 142898 344132 142986
rect 344240 142898 344420 142986
rect 344528 142898 344708 142986
rect 344816 142898 344996 142986
rect 345104 142898 345284 142986
rect 345392 142898 345572 142986
rect 345680 142898 345860 142986
rect 346114 142898 346294 142986
rect 346402 142898 346582 142986
rect 346690 142898 346870 142986
rect 346978 142898 347158 142986
rect 347266 142898 347446 142986
rect 347554 142898 347734 142986
rect 347842 142898 348022 142986
rect 348130 142898 348310 142986
rect 348564 142898 348744 142986
rect 348852 142898 349032 142986
rect 349140 142898 349320 142986
rect 349428 142898 349608 142986
rect 349716 142898 349896 142986
rect 350004 142898 350184 142986
rect 350292 142898 350472 142986
rect 350580 142898 350760 142986
rect 351014 142898 351194 142986
rect 351302 142898 351482 142986
rect 351590 142898 351770 142986
rect 351878 142898 352058 142986
rect 352166 142898 352346 142986
rect 352454 142898 352634 142986
rect 352742 142898 352922 142986
rect 353030 142898 353210 142986
rect 353464 142898 353644 142986
rect 353752 142898 353932 142986
rect 354040 142898 354220 142986
rect 354328 142898 354508 142986
rect 354616 142898 354796 142986
rect 354904 142898 355084 142986
rect 355192 142898 355372 142986
rect 355480 142898 355660 142986
rect 355914 142898 356094 142986
rect 356202 142898 356382 142986
rect 356490 142898 356670 142986
rect 356778 142898 356958 142986
rect 357066 142898 357246 142986
rect 357354 142898 357534 142986
rect 357642 142898 357822 142986
rect 357930 142898 358110 142986
rect 358364 142898 358544 142986
rect 358652 142898 358832 142986
rect 358940 142898 359120 142986
rect 359228 142898 359408 142986
rect 359516 142898 359696 142986
rect 359804 142898 359984 142986
rect 360092 142898 360272 142986
rect 360380 142898 360560 142986
rect 360814 142898 360994 142986
rect 361102 142898 361282 142986
rect 361390 142898 361570 142986
rect 361678 142898 361858 142986
rect 361966 142898 362146 142986
rect 362254 142898 362434 142986
rect 362542 142898 362722 142986
rect 362830 142898 363010 142986
rect 363264 142898 363444 142986
rect 363552 142898 363732 142986
rect 363840 142898 364020 142986
rect 364128 142898 364308 142986
rect 364416 142898 364596 142986
rect 364704 142898 364884 142986
rect 364992 142898 365172 142986
rect 365280 142898 365460 142986
rect 365714 142898 365894 142986
rect 366002 142898 366182 142986
rect 366290 142898 366470 142986
rect 366578 142898 366758 142986
rect 366866 142898 367046 142986
rect 367154 142898 367334 142986
rect 367442 142898 367622 142986
rect 367730 142898 367910 142986
<< dnwell >>
rect 242650 142250 368550 297550
<< nwell >>
rect 242550 297300 368650 297650
rect 242550 142500 242900 297300
rect 368300 142500 368650 297300
rect 242550 142150 368650 142500
<< nsubdiff >>
rect 242650 297550 242750 297575
rect 368450 297550 368550 297575
rect 242625 297450 242750 297550
rect 368450 297450 368575 297550
rect 242650 297400 242750 297450
rect 242650 142350 242750 142400
rect 368450 297400 368550 297450
rect 368450 142350 368550 142400
rect 242625 142250 242750 142350
rect 368450 142250 368575 142350
rect 242650 142225 242750 142250
rect 368450 142225 368550 142250
<< nsubdiffcont >>
rect 242750 297450 368450 297550
rect 242650 142400 242750 297400
rect 368450 142400 368550 297400
rect 242750 142250 368450 142350
<< locali >>
rect 242600 297550 368600 297600
rect 242600 297450 242750 297550
rect 368450 297450 368600 297550
rect 242600 297400 368600 297450
rect 242600 142400 242650 297400
rect 242750 142400 242800 297400
rect 368400 142400 368450 297400
rect 368550 142400 368600 297400
rect 242600 142350 368600 142400
rect 242600 142250 242750 142350
rect 368450 142250 368600 142350
rect 242600 142200 368600 142250
<< metal2 >>
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect -800 680242 1700 685242
rect 582300 677984 584800 682984
rect -800 643842 1660 648642
rect 582340 639784 584800 644584
rect -800 633842 1660 638642
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use sonos_array_50x50x64  sonos_array_50x50x64_0
timestamp 1684786423
transform 1 0 243160 0 1 142776
box -160 -176 125116 154360
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
