magic
tech sky130A
timestamp 1686033482
<< error_s >>
rect -80 1387 1250 1530
rect -80 1381 63 1387
rect 1107 1381 1250 1387
rect -80 1337 117 1381
rect 171 1337 261 1381
rect 315 1337 405 1381
rect 459 1337 549 1381
rect 603 1337 693 1381
rect 747 1337 837 1381
rect 891 1337 981 1381
rect 1035 1337 1250 1381
rect -80 1143 63 1337
rect 1107 1143 1250 1337
rect -80 1099 117 1143
rect 171 1099 261 1143
rect 315 1099 405 1143
rect 459 1099 549 1143
rect 603 1099 693 1143
rect 747 1099 837 1143
rect 891 1099 981 1143
rect 1035 1099 1250 1143
rect -80 1035 63 1099
rect 1107 1035 1250 1099
rect -80 991 117 1035
rect 171 991 261 1035
rect 315 991 405 1035
rect 459 991 549 1035
rect 603 991 693 1035
rect 747 991 837 1035
rect 891 991 981 1035
rect 1035 991 1250 1035
rect -80 797 63 991
rect 1107 797 1250 991
rect -80 753 117 797
rect 171 753 261 797
rect 315 753 405 797
rect 459 753 549 797
rect 603 753 693 797
rect 747 753 837 797
rect 891 753 981 797
rect 1035 753 1250 797
rect -80 689 63 753
rect 1107 689 1250 753
rect -80 645 117 689
rect 171 645 261 689
rect 315 645 405 689
rect 459 645 549 689
rect 603 645 693 689
rect 747 645 837 689
rect 891 645 981 689
rect 1035 645 1250 689
rect -80 451 63 645
rect 1107 451 1250 645
rect -80 407 117 451
rect 171 407 261 451
rect 315 407 405 451
rect 459 407 549 451
rect 603 407 693 451
rect 747 407 837 451
rect 891 407 981 451
rect 1035 407 1250 451
rect -80 343 63 407
rect 1107 343 1250 407
rect -80 299 117 343
rect 171 299 261 343
rect 315 299 405 343
rect 459 299 549 343
rect 603 299 693 343
rect 747 299 837 343
rect 891 299 981 343
rect 1035 299 1250 343
rect -80 105 63 299
rect 1107 105 1250 299
rect -80 61 117 105
rect 171 61 261 105
rect 315 61 405 105
rect 459 61 549 105
rect 603 61 693 105
rect 747 61 837 105
rect 891 61 981 105
rect 1035 61 1250 105
rect -80 55 63 61
rect 1107 55 1250 61
rect -80 -88 1250 55
<< dnwell >>
rect -40 -48 1210 1490
use sonos_8x8  sonos_8x8_0
timestamp 1686033482
transform 1 0 0 0 1 0
box -80 -88 1308 1530
<< end >>
