magic
tech sky130A
timestamp 1663459791
<< error_p >>
rect -42 37 42 265
rect -39 9 -16 15
rect 16 9 39 15
rect -39 -8 -36 9
rect 16 -8 19 9
rect -39 -14 -16 -8
rect 16 -14 39 -8
rect 42 -35 258 37
<< dnwell >>
rect -42 -35 42 37
<< nsonos >>
rect -42 -35 42 37
<< ndiff >>
rect -42 9 -11 23
rect -42 -8 -36 9
rect -19 -8 -11 9
rect -42 -22 -11 -8
rect 11 9 42 23
rect 11 -8 19 9
rect 36 -8 42 9
rect 11 -22 42 -8
<< ndiffc >>
rect -36 -8 -19 9
rect 19 -8 36 9
<< poly >>
rect -11 23 11 37
rect -11 -35 11 -22
<< locali >>
rect -36 9 -19 17
rect -36 -16 -19 -8
rect 19 9 36 17
rect 19 -16 36 -8
<< viali >>
rect -36 -8 -19 9
rect 19 -8 36 9
<< metal1 >>
rect -39 9 -16 15
rect -39 -8 -36 9
rect -19 -8 -16 9
rect -39 -14 -16 -8
rect 16 9 39 15
rect 16 -8 19 9
rect 36 -8 39 9
rect 16 -14 39 -8
<< properties >>
string FIXED_BBOX -84 -70 84 70
string gencell sky130_fd_bs_flash__special_sonosfet_star
string library sky130
string parameters w 0.450 l 0.22 m 1 nf 1 diffcov 50 polycov 50 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 50 viadrn 50 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
