magic
tech sky130A
magscale 1 2
timestamp 1663041771
<< error_s >>
rect -249 1341 1401 1467
rect -249 -339 -123 1341
rect 27 1052 117 1096
rect 171 1052 261 1096
rect 315 1052 405 1096
rect 459 1052 549 1096
rect 603 1052 693 1096
rect 747 1052 837 1096
rect 891 1052 981 1096
rect 1035 1052 1125 1096
rect 27 944 117 988
rect 171 944 261 988
rect 315 944 405 988
rect 459 944 549 988
rect 603 944 693 988
rect 747 944 837 988
rect 891 944 981 988
rect 1035 944 1125 988
rect 27 706 117 750
rect 171 706 261 750
rect 315 706 405 750
rect 459 706 549 750
rect 603 706 693 750
rect 747 706 837 750
rect 891 706 981 750
rect 1035 706 1125 750
rect 27 598 117 642
rect 171 598 261 642
rect 315 598 405 642
rect 459 598 549 642
rect 603 598 693 642
rect 747 598 837 642
rect 891 598 981 642
rect 1035 598 1125 642
rect 27 360 117 404
rect 171 360 261 404
rect 315 360 405 404
rect 459 360 549 404
rect 603 360 693 404
rect 747 360 837 404
rect 891 360 981 404
rect 1035 360 1125 404
rect 27 252 117 296
rect 171 252 261 296
rect 315 252 405 296
rect 459 252 549 296
rect 603 252 693 296
rect 747 252 837 296
rect 891 252 981 296
rect 1035 252 1125 296
rect 27 14 117 58
rect 171 14 261 58
rect 315 14 405 58
rect 459 14 549 58
rect 603 14 693 58
rect 747 14 837 58
rect 891 14 981 58
rect 1035 14 1125 58
rect 27 -94 117 -50
rect 171 -94 261 -50
rect 315 -94 405 -50
rect 459 -94 549 -50
rect 603 -94 693 -50
rect 747 -94 837 -50
rect 891 -94 981 -50
rect 1035 -94 1125 -50
rect 1275 -339 1401 1341
rect -249 -465 1401 -339
<< dnwell >>
rect 0 -32 1 177
<< poly >>
rect 0 100 1 130
rect 0 14 1 58
use sonos_array_corner  sonos_array_corner_0
timestamp 1663041771
transform 1 0 0 0 1 0
box -417 -633 271 55
use sonos_array_corner  sonos_array_corner_1
timestamp 1663041771
transform 1 0 0 0 -1 1002
box -417 -633 271 55
use sonos_array_corner  sonos_array_corner_2
timestamp 1663041771
transform -1 0 1152 0 1 0
box -417 -633 271 55
use sonos_array_corner  sonos_array_corner_3
timestamp 1663041771
transform -1 0 1152 0 -1 1002
box -417 -633 271 55
use sonos_cell  sonos_cell_0
array 0 7 144 0 3 346
timestamp 1663041771
transform 1 0 72 0 1 79
box -152 -206 528 474
use sonos_cell  sonos_cell_1
array 0 7 144 0 3 -346
timestamp 1663041771
transform 1 0 72 0 -1 -115
box -152 -206 528 474
use sonos_endcap_lr  sonos_endcap_lr_0
array 0 0 417 0 3 346
timestamp 1663041771
transform 1 0 0 0 1 0
box -417 -292 271 388
use sonos_endcap_lr  sonos_endcap_lr_1
array 0 0 417 0 3 346
timestamp 1663041771
transform -1 0 1152 0 -1 1002
box -417 -292 271 388
use sonos_endcap_tb  sonos_endcap_tb_0
array 0 7 144 0 0 154
timestamp 1663041771
transform 1 0 204 0 1 215
box -284 -848 396 -160
use sonos_endcap_tb  sonos_endcap_tb_1
array 0 7 144 0 0 -154
timestamp 1663041771
transform 1 0 204 0 -1 787
box -284 -848 396 -160
<< labels >>
rlabel space -417 -187 -381 -153 1 wl0
rlabel space -417 -113 -381 -79 1 wls0
rlabel space 1533 -93 1569 -59 1 wls0
rlabel space 1533 -161 1569 -127 1 nc0
rlabel space -417 -45 -381 -11 1 nc0
rlabel space -417 23 -381 57 1 wls1
rlabel space 1533 43 1569 77 1 wls1
rlabel space 1533 -25 1569 9 1 nc1
rlabel space -417 91 -381 125 1 nc1
rlabel space 1533 185 1569 219 1 nc2
rlabel space 1533 117 1569 151 1 wl1
rlabel space -417 159 -381 193 1 wl2
rlabel space -417 233 -381 267 1 wls2
rlabel space 1533 253 1569 287 1 wls2
rlabel space 1533 321 1569 355 1 nc3
rlabel space -417 301 -381 335 1 nc2
rlabel space -417 369 -381 403 1 wls3
rlabel space -417 437 -381 471 1 nc3
rlabel space -417 505 -381 539 1 wl4
rlabel space 1533 389 1569 423 1 wls3
rlabel space 1533 463 1569 497 1 wl3
rlabel space 1533 531 1569 565 1 nc4
rlabel space 1533 667 1569 701 1 nc5
rlabel space 1533 877 1569 911 1 nc6
rlabel space 1533 1013 1569 1047 1 nc7
rlabel space 1533 599 1569 633 1 wls4
rlabel space -417 579 -381 613 1 wls4
rlabel space -417 647 -381 681 1 nc4
rlabel space -417 783 -381 817 1 nc5
rlabel space -417 993 -381 1027 1 nc6
rlabel space -417 1129 -381 1163 1 nc7
rlabel space 1533 735 1569 769 1 wls5
rlabel space -417 715 -381 749 1 wls5
rlabel space 1533 809 1569 843 1 wl5
rlabel space -417 851 -381 885 1 wl6
rlabel space 1533 945 1569 979 1 wls6
rlabel space -417 925 -381 959 1 wls6
rlabel space -417 1061 -381 1095 1 wls7
rlabel space 1533 1081 1569 1115 1 wls7
rlabel space 1533 1155 1569 1189 1 wl7
rlabel space 54 -633 90 -597 1 bl0
rlabel space 124 -633 160 -597 1 src0
rlabel space 198 -633 234 -597 1 bl1
rlabel space 268 -633 304 -597 1 src1
rlabel space 342 -633 378 -597 1 bl2
rlabel space 412 -633 448 -597 1 src2
rlabel space 486 -633 522 -597 1 bl3
rlabel space 556 -633 592 -597 1 src3
rlabel space 630 -633 666 -597 1 bl4
rlabel space 700 -633 736 -597 1 src4
rlabel space 774 -633 810 -597 1 bl5
rlabel space 844 -633 880 -597 1 src5
rlabel space 918 -633 954 -597 1 bl6
rlabel space 988 -633 1024 -597 1 src6
rlabel space 1062 -633 1098 -597 1 bl7
rlabel space 1132 -633 1168 -597 1 src7
rlabel space 54 1599 90 1635 1 bl0
rlabel space 124 1599 160 1635 1 src0
rlabel space 198 1599 234 1635 1 bl1
rlabel space 268 1599 304 1635 1 src1
rlabel space 342 1599 378 1635 1 bl2
rlabel space 412 1599 448 1635 1 src2
rlabel space 486 1599 522 1635 1 bl3
rlabel space 556 1599 592 1635 1 src3
rlabel space 630 1599 666 1635 1 bl4
rlabel space 700 1599 736 1635 1 src4
rlabel space 774 1599 810 1635 1 bl5
rlabel space 844 1599 880 1635 1 src5
rlabel space 918 1599 954 1635 1 bl6
rlabel space 988 1599 1024 1635 1 src6
rlabel space 1062 1599 1098 1635 1 bl7
rlabel space 1132 1599 1168 1635 1 src7
rlabel space -111 1382 -50 1440 1 B
rlabel space 1202 1382 1263 1440 1 B
rlabel space 1202 -438 1263 -380 1 B
rlabel space -111 -439 -50 -381 1 B
<< end >>
