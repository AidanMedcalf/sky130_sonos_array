magic
tech sky130A
timestamp 1663090256
<< checkpaint >>
rect -284 -979 396 -293
<< dnwell >>
rect -204 -893 -59 -680
rect -204 -680 -60 -373
<< nwell >>
rect -204 -979 -60 -680
<< nsubdiff >>
rect -204 -943 -60 -938
rect -204 -938 -187 -904
rect -77 -938 -60 -904
rect -204 -904 -60 -898
<< nsubdiffcont >>
rect -187 -938 -77 -904
<< locali >>
rect -204 -938 -187 -904
rect -77 -938 -60 -904
rect -204 -629 -149 -595
rect -115 -629 -59 -595
rect -154 -519 -111 -503
rect -154 -503 -149 -469
rect -115 -503 -111 -469
rect -154 -469 -111 -439
rect -154 -439 -44 -423
rect -154 -423 -149 -389
rect -115 -423 -79 -389
rect -45 -423 -44 -389
rect -154 -389 -44 -373
<< viali >>
rect -79 -423 -45 -389
<< metal1 >>
rect -150 -943 -114 -381
rect -80 -943 -44 -429
rect -85 -429 -39 -423
rect -85 -423 -79 -389
rect -45 -423 -39 -389
rect -85 -389 -39 -383
rect -80 -383 -44 -377
<< poly >>
rect -204 -461 -177 -431
rect -87 -461 -60 -431
<< error_p >>
rect -240 -979 -204 -973
rect -60 -979 -24 -973
rect -284 -973 -204 -943
rect -187 -962 -163 -943
rect -101 -962 -77 -943
rect -60 -973 21 -943
rect -284 -943 -168 -898
rect -96 -943 21 -898
rect -60 -898 21 -893
rect -187 -898 -163 -880
rect -101 -898 -77 -880
rect -284 -898 -204 -680
rect -60 -893 396 -680
rect -284 -680 396 -373
rect -284 -373 20 -293
<< psubdiff >>
rect -204 -653 -59 -629
rect -204 -629 -149 -595
rect -115 -629 -59 -595
rect -204 -595 -59 -577
<< ndiff >>
rect -177 -523 -87 -503
rect -177 -503 -149 -469
rect -115 -503 -87 -469
rect -177 -469 -87 -461
rect -177 -431 -87 -423
rect -177 -423 -149 -389
rect -115 -423 -87 -389
rect -177 -389 -87 -381
<< ndiffc >>
rect -149 -503 -115 -469
rect -149 -423 -115 -389
<< psubdiffcont >>
rect -149 -629 -115 -595
<< npd >>
rect -177 -461 -87 -431
<< end >>
