magic
tech sky130A
timestamp 1685567320
<< dnwell >>
rect -2 0 514 522
<< nwell >>
rect -57 419 569 577
rect -57 103 101 419
rect 411 103 569 419
rect -57 -55 569 103
<< pwell >>
rect -100 577 612 620
rect -100 -55 -57 577
rect 569 -55 612 577
rect -100 -98 612 -55
<< mvpsubdiff >>
rect -118 620 17 638
rect 495 620 630 638
rect -118 503 -100 620
rect -118 -98 -100 19
rect 612 503 630 620
rect 612 -98 630 19
rect -118 -116 17 -98
rect 495 -116 630 -98
<< mvnsubdiff >>
rect -24 534 536 544
rect -24 516 17 534
rect 495 516 536 534
rect -24 506 536 516
rect -24 503 14 506
rect -24 19 -14 503
rect 4 19 14 503
rect -24 16 14 19
rect 498 503 536 506
rect 498 19 508 503
rect 526 19 536 503
rect 498 16 536 19
rect -24 6 536 16
rect -24 -12 17 6
rect 495 -12 536 6
rect -24 -22 536 -12
<< mvpsubdiffcont >>
rect 17 620 495 638
rect -118 19 -100 503
rect 612 19 630 503
rect 17 -116 495 -98
<< mvnsubdiffcont >>
rect 17 516 495 534
rect -14 19 4 503
rect 508 19 526 503
rect 17 -12 495 6
<< locali >>
rect -118 620 17 638
rect 495 620 630 638
rect -118 503 -100 620
rect -118 -98 -100 19
rect -14 516 17 534
rect 495 516 526 534
rect -14 503 4 516
rect -14 6 4 19
rect 508 503 526 516
rect 508 6 526 19
rect -14 -12 17 6
rect 495 -12 526 6
rect 612 503 630 620
rect 612 -98 630 19
rect -118 -116 17 -98
rect 495 -116 630 -98
<< metal1 >>
rect 238 283 274 308
use sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_bs_flash__special_sonosfet_star_0
timestamp 1685564080
transform 1 0 256 0 1 261
box -258 -261 258 261
<< labels >>
flabel metal1 238 283 274 308 1 FreeSans 144 0 0 -64 G
flabel metal1 220 239 237 253 1 FreeSans 144 0 0 -80 S
flabel metal1 275 239 292 253 1 FreeSans 144 0 0 -80 D
flabel locali -14 520 4 534 1 FreeSans 144 0 0 -80 VNB
flabel locali 165 341 182 355 1 FreeSans 144 0 0 -80 B
flabel locali -118 624 -100 638 1 FreeSans 144 0 0 -80 VPB
<< properties >>
string FIXED_BBOX -5 517 -4 525
<< end >>
