magic
tech sky130A
magscale 1 2
timestamp 1663041771
<< error_s >>
rect 168 1974 1818 2100
rect 168 294 294 1974
rect 444 1685 534 1729
rect 588 1685 678 1729
rect 732 1685 822 1729
rect 876 1685 966 1729
rect 1020 1685 1110 1729
rect 1164 1685 1254 1729
rect 1308 1685 1398 1729
rect 1452 1685 1542 1729
rect 444 1577 534 1621
rect 588 1577 678 1621
rect 732 1577 822 1621
rect 876 1577 966 1621
rect 1020 1577 1110 1621
rect 1164 1577 1254 1621
rect 1308 1577 1398 1621
rect 1452 1577 1542 1621
rect 444 1339 534 1383
rect 588 1339 678 1383
rect 732 1339 822 1383
rect 876 1339 966 1383
rect 1020 1339 1110 1383
rect 1164 1339 1254 1383
rect 1308 1339 1398 1383
rect 1452 1339 1542 1383
rect 444 1231 534 1275
rect 588 1231 678 1275
rect 732 1231 822 1275
rect 876 1231 966 1275
rect 1020 1231 1110 1275
rect 1164 1231 1254 1275
rect 1308 1231 1398 1275
rect 1452 1231 1542 1275
rect 444 993 534 1037
rect 588 993 678 1037
rect 732 993 822 1037
rect 876 993 966 1037
rect 1020 993 1110 1037
rect 1164 993 1254 1037
rect 1308 993 1398 1037
rect 1452 993 1542 1037
rect 444 885 534 929
rect 588 885 678 929
rect 732 885 822 929
rect 876 885 966 929
rect 1020 885 1110 929
rect 1164 885 1254 929
rect 1308 885 1398 929
rect 1452 885 1542 929
rect 444 647 534 691
rect 588 647 678 691
rect 732 647 822 691
rect 876 647 966 691
rect 1020 647 1110 691
rect 1164 647 1254 691
rect 1308 647 1398 691
rect 1452 647 1542 691
rect 444 539 534 583
rect 588 539 678 583
rect 732 539 822 583
rect 876 539 966 583
rect 1020 539 1110 583
rect 1164 539 1254 583
rect 1308 539 1398 583
rect 1452 539 1542 583
rect 1692 294 1818 1974
rect 168 168 1818 294
<< metal1 >>
rect 464 2290 1592 2296
rect 464 2238 470 2290
rect 1586 2238 1592 2290
rect 464 2232 1592 2238
rect 1950 1822 2014 1828
rect -28 1796 36 1802
rect -28 438 -22 1796
rect 30 438 36 1796
rect 1950 472 1956 1822
rect 2008 472 2014 1822
rect 1950 466 2014 472
rect -28 432 36 438
rect 464 30 1592 36
rect 464 -22 470 30
rect 1586 -22 1592 30
rect 464 -28 1592 -22
<< via1 >>
rect 470 2238 1586 2290
rect -22 438 30 1796
rect 1956 472 2008 1822
rect 470 -22 1586 30
<< metal2 >>
rect -30 2290 2014 2296
rect -30 2238 470 2290
rect 1586 2238 2014 2290
rect -30 1822 2014 2238
rect -30 1796 1956 1822
rect -30 438 -22 1796
rect 30 472 1956 1796
rect 2008 472 2014 1822
rect 30 438 2014 472
rect -30 30 2014 438
rect -30 -22 470 30
rect 1586 -22 2014 30
rect -30 -28 2014 -22
use sonos_array  sonos_array_0
timestamp 1663041771
transform 1 0 417 0 1 633
box -417 -633 1608 1635
<< labels >>
rlabel metal2 -30 -28 2014 2296 1 vss
<< end >>
