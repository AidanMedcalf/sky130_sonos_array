magic
tech sky130A
timestamp 1663354744
<< metal1 >>
rect 0 412 165 458
rect 54 404 90 412
rect 124 400 160 412
<< end >>
