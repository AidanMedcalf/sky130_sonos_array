magic
tech sky130A
timestamp 1663450679
<< error_p >>
rect -40 1442 1192 1482
rect -40 0 1308 1442
rect -40 -40 1192 0
use sonos_cell_mirrored  sonos_cell_mirrored_0
array 0 7 144 0 3 346
timestamp 1663450679
transform 1 0 -80 0 1 -80
box 40 40 380 524
<< end >>
