magic
tech sky130A
magscale 1 2
timestamp 1685138211
<< error_p >>
rect 180350 326988 180530 327076
rect 180638 326988 180818 327076
rect 180926 326988 181106 327076
rect 181214 326988 181394 327076
rect 181502 326988 181682 327076
rect 181790 326988 181970 327076
rect 182078 326988 182258 327076
rect 182366 326988 182546 327076
rect 194846 326988 195026 327076
rect 195134 326988 195314 327076
rect 195422 326988 195602 327076
rect 195710 326988 195890 327076
rect 195998 326988 196178 327076
rect 196286 326988 196466 327076
rect 196574 326988 196754 327076
rect 196862 326988 197042 327076
rect 209342 326988 209522 327076
rect 209630 326988 209810 327076
rect 209918 326988 210098 327076
rect 210206 326988 210386 327076
rect 210494 326988 210674 327076
rect 210782 326988 210962 327076
rect 211070 326988 211250 327076
rect 211358 326988 211538 327076
rect 223838 326988 224018 327076
rect 224126 326988 224306 327076
rect 224414 326988 224594 327076
rect 224702 326988 224882 327076
rect 224990 326988 225170 327076
rect 225278 326988 225458 327076
rect 225566 326988 225746 327076
rect 225854 326988 226034 327076
rect 238334 326988 238514 327076
rect 238622 326988 238802 327076
rect 238910 326988 239090 327076
rect 239198 326988 239378 327076
rect 239486 326988 239666 327076
rect 239774 326988 239954 327076
rect 240062 326988 240242 327076
rect 240350 326988 240530 327076
rect 252830 326988 253010 327076
rect 253118 326988 253298 327076
rect 253406 326988 253586 327076
rect 253694 326988 253874 327076
rect 253982 326988 254162 327076
rect 254270 326988 254450 327076
rect 254558 326988 254738 327076
rect 254846 326988 255026 327076
rect 267326 326988 267506 327076
rect 267614 326988 267794 327076
rect 267902 326988 268082 327076
rect 268190 326988 268370 327076
rect 268478 326988 268658 327076
rect 268766 326988 268946 327076
rect 269054 326988 269234 327076
rect 269342 326988 269522 327076
rect 281822 326988 282002 327076
rect 282110 326988 282290 327076
rect 282398 326988 282578 327076
rect 282686 326988 282866 327076
rect 282974 326988 283154 327076
rect 283262 326988 283442 327076
rect 283550 326988 283730 327076
rect 283838 326988 284018 327076
rect 296318 326988 296498 327076
rect 296606 326988 296786 327076
rect 296894 326988 297074 327076
rect 297182 326988 297362 327076
rect 297470 326988 297650 327076
rect 297758 326988 297938 327076
rect 298046 326988 298226 327076
rect 298334 326988 298514 327076
rect 310814 326988 310994 327076
rect 311102 326988 311282 327076
rect 311390 326988 311570 327076
rect 311678 326988 311858 327076
rect 311966 326988 312146 327076
rect 312254 326988 312434 327076
rect 312542 326988 312722 327076
rect 312830 326988 313010 327076
rect 325310 326988 325490 327076
rect 325598 326988 325778 327076
rect 325886 326988 326066 327076
rect 326174 326988 326354 327076
rect 326462 326988 326642 327076
rect 326750 326988 326930 327076
rect 327038 326988 327218 327076
rect 327326 326988 327506 327076
rect 339806 326988 339986 327076
rect 340094 326988 340274 327076
rect 340382 326988 340562 327076
rect 340670 326988 340850 327076
rect 340958 326988 341138 327076
rect 341246 326988 341426 327076
rect 341534 326988 341714 327076
rect 341822 326988 342002 327076
rect 354302 326988 354482 327076
rect 354590 326988 354770 327076
rect 354878 326988 355058 327076
rect 355166 326988 355346 327076
rect 355454 326988 355634 327076
rect 355742 326988 355922 327076
rect 356030 326988 356210 327076
rect 356318 326988 356498 327076
rect 368798 326988 368978 327076
rect 369086 326988 369266 327076
rect 369374 326988 369554 327076
rect 369662 326988 369842 327076
rect 369950 326988 370130 327076
rect 370238 326988 370418 327076
rect 370526 326988 370706 327076
rect 370814 326988 370994 327076
rect 383294 326988 383474 327076
rect 383582 326988 383762 327076
rect 383870 326988 384050 327076
rect 384158 326988 384338 327076
rect 384446 326988 384626 327076
rect 384734 326988 384914 327076
rect 385022 326988 385202 327076
rect 385310 326988 385490 327076
rect 397790 326988 397970 327076
rect 398078 326988 398258 327076
rect 398366 326988 398546 327076
rect 398654 326988 398834 327076
rect 398942 326988 399122 327076
rect 399230 326988 399410 327076
rect 399518 326988 399698 327076
rect 399806 326988 399986 327076
rect 412286 326988 412466 327076
rect 412574 326988 412754 327076
rect 412862 326988 413042 327076
rect 413150 326988 413330 327076
rect 413438 326988 413618 327076
rect 413726 326988 413906 327076
rect 414014 326988 414194 327076
rect 414302 326988 414482 327076
rect 426782 326988 426962 327076
rect 427070 326988 427250 327076
rect 427358 326988 427538 327076
rect 427646 326988 427826 327076
rect 427934 326988 428114 327076
rect 428222 326988 428402 327076
rect 428510 326988 428690 327076
rect 428798 326988 428978 327076
rect 441278 326988 441458 327076
rect 441566 326988 441746 327076
rect 441854 326988 442034 327076
rect 442142 326988 442322 327076
rect 442430 326988 442610 327076
rect 442718 326988 442898 327076
rect 443006 326988 443186 327076
rect 443294 326988 443474 327076
rect 455774 326988 455954 327076
rect 456062 326988 456242 327076
rect 456350 326988 456530 327076
rect 456638 326988 456818 327076
rect 456926 326988 457106 327076
rect 457214 326988 457394 327076
rect 457502 326988 457682 327076
rect 457790 326988 457970 327076
rect 180350 326772 180530 326860
rect 180638 326772 180818 326860
rect 180926 326772 181106 326860
rect 181214 326772 181394 326860
rect 181502 326772 181682 326860
rect 181790 326772 181970 326860
rect 182078 326772 182258 326860
rect 182366 326772 182546 326860
rect 194846 326772 195026 326860
rect 195134 326772 195314 326860
rect 195422 326772 195602 326860
rect 195710 326772 195890 326860
rect 195998 326772 196178 326860
rect 196286 326772 196466 326860
rect 196574 326772 196754 326860
rect 196862 326772 197042 326860
rect 209342 326772 209522 326860
rect 209630 326772 209810 326860
rect 209918 326772 210098 326860
rect 210206 326772 210386 326860
rect 210494 326772 210674 326860
rect 210782 326772 210962 326860
rect 211070 326772 211250 326860
rect 211358 326772 211538 326860
rect 223838 326772 224018 326860
rect 224126 326772 224306 326860
rect 224414 326772 224594 326860
rect 224702 326772 224882 326860
rect 224990 326772 225170 326860
rect 225278 326772 225458 326860
rect 225566 326772 225746 326860
rect 225854 326772 226034 326860
rect 238334 326772 238514 326860
rect 238622 326772 238802 326860
rect 238910 326772 239090 326860
rect 239198 326772 239378 326860
rect 239486 326772 239666 326860
rect 239774 326772 239954 326860
rect 240062 326772 240242 326860
rect 240350 326772 240530 326860
rect 252830 326772 253010 326860
rect 253118 326772 253298 326860
rect 253406 326772 253586 326860
rect 253694 326772 253874 326860
rect 253982 326772 254162 326860
rect 254270 326772 254450 326860
rect 254558 326772 254738 326860
rect 254846 326772 255026 326860
rect 267326 326772 267506 326860
rect 267614 326772 267794 326860
rect 267902 326772 268082 326860
rect 268190 326772 268370 326860
rect 268478 326772 268658 326860
rect 268766 326772 268946 326860
rect 269054 326772 269234 326860
rect 269342 326772 269522 326860
rect 281822 326772 282002 326860
rect 282110 326772 282290 326860
rect 282398 326772 282578 326860
rect 282686 326772 282866 326860
rect 282974 326772 283154 326860
rect 283262 326772 283442 326860
rect 283550 326772 283730 326860
rect 283838 326772 284018 326860
rect 296318 326772 296498 326860
rect 296606 326772 296786 326860
rect 296894 326772 297074 326860
rect 297182 326772 297362 326860
rect 297470 326772 297650 326860
rect 297758 326772 297938 326860
rect 298046 326772 298226 326860
rect 298334 326772 298514 326860
rect 310814 326772 310994 326860
rect 311102 326772 311282 326860
rect 311390 326772 311570 326860
rect 311678 326772 311858 326860
rect 311966 326772 312146 326860
rect 312254 326772 312434 326860
rect 312542 326772 312722 326860
rect 312830 326772 313010 326860
rect 325310 326772 325490 326860
rect 325598 326772 325778 326860
rect 325886 326772 326066 326860
rect 326174 326772 326354 326860
rect 326462 326772 326642 326860
rect 326750 326772 326930 326860
rect 327038 326772 327218 326860
rect 327326 326772 327506 326860
rect 339806 326772 339986 326860
rect 340094 326772 340274 326860
rect 340382 326772 340562 326860
rect 340670 326772 340850 326860
rect 340958 326772 341138 326860
rect 341246 326772 341426 326860
rect 341534 326772 341714 326860
rect 341822 326772 342002 326860
rect 354302 326772 354482 326860
rect 354590 326772 354770 326860
rect 354878 326772 355058 326860
rect 355166 326772 355346 326860
rect 355454 326772 355634 326860
rect 355742 326772 355922 326860
rect 356030 326772 356210 326860
rect 356318 326772 356498 326860
rect 368798 326772 368978 326860
rect 369086 326772 369266 326860
rect 369374 326772 369554 326860
rect 369662 326772 369842 326860
rect 369950 326772 370130 326860
rect 370238 326772 370418 326860
rect 370526 326772 370706 326860
rect 370814 326772 370994 326860
rect 383294 326772 383474 326860
rect 383582 326772 383762 326860
rect 383870 326772 384050 326860
rect 384158 326772 384338 326860
rect 384446 326772 384626 326860
rect 384734 326772 384914 326860
rect 385022 326772 385202 326860
rect 385310 326772 385490 326860
rect 397790 326772 397970 326860
rect 398078 326772 398258 326860
rect 398366 326772 398546 326860
rect 398654 326772 398834 326860
rect 398942 326772 399122 326860
rect 399230 326772 399410 326860
rect 399518 326772 399698 326860
rect 399806 326772 399986 326860
rect 412286 326772 412466 326860
rect 412574 326772 412754 326860
rect 412862 326772 413042 326860
rect 413150 326772 413330 326860
rect 413438 326772 413618 326860
rect 413726 326772 413906 326860
rect 414014 326772 414194 326860
rect 414302 326772 414482 326860
rect 426782 326772 426962 326860
rect 427070 326772 427250 326860
rect 427358 326772 427538 326860
rect 427646 326772 427826 326860
rect 427934 326772 428114 326860
rect 428222 326772 428402 326860
rect 428510 326772 428690 326860
rect 428798 326772 428978 326860
rect 441278 326772 441458 326860
rect 441566 326772 441746 326860
rect 441854 326772 442034 326860
rect 442142 326772 442322 326860
rect 442430 326772 442610 326860
rect 442718 326772 442898 326860
rect 443006 326772 443186 326860
rect 443294 326772 443474 326860
rect 455774 326772 455954 326860
rect 456062 326772 456242 326860
rect 456350 326772 456530 326860
rect 456638 326772 456818 326860
rect 456926 326772 457106 326860
rect 457214 326772 457394 326860
rect 457502 326772 457682 326860
rect 457790 326772 457970 326860
rect 180350 326296 180530 326384
rect 180638 326296 180818 326384
rect 180926 326296 181106 326384
rect 181214 326296 181394 326384
rect 181502 326296 181682 326384
rect 181790 326296 181970 326384
rect 182078 326296 182258 326384
rect 182366 326296 182546 326384
rect 194846 326296 195026 326384
rect 195134 326296 195314 326384
rect 195422 326296 195602 326384
rect 195710 326296 195890 326384
rect 195998 326296 196178 326384
rect 196286 326296 196466 326384
rect 196574 326296 196754 326384
rect 196862 326296 197042 326384
rect 209342 326296 209522 326384
rect 209630 326296 209810 326384
rect 209918 326296 210098 326384
rect 210206 326296 210386 326384
rect 210494 326296 210674 326384
rect 210782 326296 210962 326384
rect 211070 326296 211250 326384
rect 211358 326296 211538 326384
rect 223838 326296 224018 326384
rect 224126 326296 224306 326384
rect 224414 326296 224594 326384
rect 224702 326296 224882 326384
rect 224990 326296 225170 326384
rect 225278 326296 225458 326384
rect 225566 326296 225746 326384
rect 225854 326296 226034 326384
rect 238334 326296 238514 326384
rect 238622 326296 238802 326384
rect 238910 326296 239090 326384
rect 239198 326296 239378 326384
rect 239486 326296 239666 326384
rect 239774 326296 239954 326384
rect 240062 326296 240242 326384
rect 240350 326296 240530 326384
rect 252830 326296 253010 326384
rect 253118 326296 253298 326384
rect 253406 326296 253586 326384
rect 253694 326296 253874 326384
rect 253982 326296 254162 326384
rect 254270 326296 254450 326384
rect 254558 326296 254738 326384
rect 254846 326296 255026 326384
rect 267326 326296 267506 326384
rect 267614 326296 267794 326384
rect 267902 326296 268082 326384
rect 268190 326296 268370 326384
rect 268478 326296 268658 326384
rect 268766 326296 268946 326384
rect 269054 326296 269234 326384
rect 269342 326296 269522 326384
rect 281822 326296 282002 326384
rect 282110 326296 282290 326384
rect 282398 326296 282578 326384
rect 282686 326296 282866 326384
rect 282974 326296 283154 326384
rect 283262 326296 283442 326384
rect 283550 326296 283730 326384
rect 283838 326296 284018 326384
rect 296318 326296 296498 326384
rect 296606 326296 296786 326384
rect 296894 326296 297074 326384
rect 297182 326296 297362 326384
rect 297470 326296 297650 326384
rect 297758 326296 297938 326384
rect 298046 326296 298226 326384
rect 298334 326296 298514 326384
rect 310814 326296 310994 326384
rect 311102 326296 311282 326384
rect 311390 326296 311570 326384
rect 311678 326296 311858 326384
rect 311966 326296 312146 326384
rect 312254 326296 312434 326384
rect 312542 326296 312722 326384
rect 312830 326296 313010 326384
rect 325310 326296 325490 326384
rect 325598 326296 325778 326384
rect 325886 326296 326066 326384
rect 326174 326296 326354 326384
rect 326462 326296 326642 326384
rect 326750 326296 326930 326384
rect 327038 326296 327218 326384
rect 327326 326296 327506 326384
rect 339806 326296 339986 326384
rect 340094 326296 340274 326384
rect 340382 326296 340562 326384
rect 340670 326296 340850 326384
rect 340958 326296 341138 326384
rect 341246 326296 341426 326384
rect 341534 326296 341714 326384
rect 341822 326296 342002 326384
rect 354302 326296 354482 326384
rect 354590 326296 354770 326384
rect 354878 326296 355058 326384
rect 355166 326296 355346 326384
rect 355454 326296 355634 326384
rect 355742 326296 355922 326384
rect 356030 326296 356210 326384
rect 356318 326296 356498 326384
rect 368798 326296 368978 326384
rect 369086 326296 369266 326384
rect 369374 326296 369554 326384
rect 369662 326296 369842 326384
rect 369950 326296 370130 326384
rect 370238 326296 370418 326384
rect 370526 326296 370706 326384
rect 370814 326296 370994 326384
rect 383294 326296 383474 326384
rect 383582 326296 383762 326384
rect 383870 326296 384050 326384
rect 384158 326296 384338 326384
rect 384446 326296 384626 326384
rect 384734 326296 384914 326384
rect 385022 326296 385202 326384
rect 385310 326296 385490 326384
rect 397790 326296 397970 326384
rect 398078 326296 398258 326384
rect 398366 326296 398546 326384
rect 398654 326296 398834 326384
rect 398942 326296 399122 326384
rect 399230 326296 399410 326384
rect 399518 326296 399698 326384
rect 399806 326296 399986 326384
rect 412286 326296 412466 326384
rect 412574 326296 412754 326384
rect 412862 326296 413042 326384
rect 413150 326296 413330 326384
rect 413438 326296 413618 326384
rect 413726 326296 413906 326384
rect 414014 326296 414194 326384
rect 414302 326296 414482 326384
rect 426782 326296 426962 326384
rect 427070 326296 427250 326384
rect 427358 326296 427538 326384
rect 427646 326296 427826 326384
rect 427934 326296 428114 326384
rect 428222 326296 428402 326384
rect 428510 326296 428690 326384
rect 428798 326296 428978 326384
rect 441278 326296 441458 326384
rect 441566 326296 441746 326384
rect 441854 326296 442034 326384
rect 442142 326296 442322 326384
rect 442430 326296 442610 326384
rect 442718 326296 442898 326384
rect 443006 326296 443186 326384
rect 443294 326296 443474 326384
rect 455774 326296 455954 326384
rect 456062 326296 456242 326384
rect 456350 326296 456530 326384
rect 456638 326296 456818 326384
rect 456926 326296 457106 326384
rect 457214 326296 457394 326384
rect 457502 326296 457682 326384
rect 457790 326296 457970 326384
rect 180350 326080 180530 326168
rect 180638 326080 180818 326168
rect 180926 326080 181106 326168
rect 181214 326080 181394 326168
rect 181502 326080 181682 326168
rect 181790 326080 181970 326168
rect 182078 326080 182258 326168
rect 182366 326080 182546 326168
rect 194846 326080 195026 326168
rect 195134 326080 195314 326168
rect 195422 326080 195602 326168
rect 195710 326080 195890 326168
rect 195998 326080 196178 326168
rect 196286 326080 196466 326168
rect 196574 326080 196754 326168
rect 196862 326080 197042 326168
rect 209342 326080 209522 326168
rect 209630 326080 209810 326168
rect 209918 326080 210098 326168
rect 210206 326080 210386 326168
rect 210494 326080 210674 326168
rect 210782 326080 210962 326168
rect 211070 326080 211250 326168
rect 211358 326080 211538 326168
rect 223838 326080 224018 326168
rect 224126 326080 224306 326168
rect 224414 326080 224594 326168
rect 224702 326080 224882 326168
rect 224990 326080 225170 326168
rect 225278 326080 225458 326168
rect 225566 326080 225746 326168
rect 225854 326080 226034 326168
rect 238334 326080 238514 326168
rect 238622 326080 238802 326168
rect 238910 326080 239090 326168
rect 239198 326080 239378 326168
rect 239486 326080 239666 326168
rect 239774 326080 239954 326168
rect 240062 326080 240242 326168
rect 240350 326080 240530 326168
rect 252830 326080 253010 326168
rect 253118 326080 253298 326168
rect 253406 326080 253586 326168
rect 253694 326080 253874 326168
rect 253982 326080 254162 326168
rect 254270 326080 254450 326168
rect 254558 326080 254738 326168
rect 254846 326080 255026 326168
rect 267326 326080 267506 326168
rect 267614 326080 267794 326168
rect 267902 326080 268082 326168
rect 268190 326080 268370 326168
rect 268478 326080 268658 326168
rect 268766 326080 268946 326168
rect 269054 326080 269234 326168
rect 269342 326080 269522 326168
rect 281822 326080 282002 326168
rect 282110 326080 282290 326168
rect 282398 326080 282578 326168
rect 282686 326080 282866 326168
rect 282974 326080 283154 326168
rect 283262 326080 283442 326168
rect 283550 326080 283730 326168
rect 283838 326080 284018 326168
rect 296318 326080 296498 326168
rect 296606 326080 296786 326168
rect 296894 326080 297074 326168
rect 297182 326080 297362 326168
rect 297470 326080 297650 326168
rect 297758 326080 297938 326168
rect 298046 326080 298226 326168
rect 298334 326080 298514 326168
rect 310814 326080 310994 326168
rect 311102 326080 311282 326168
rect 311390 326080 311570 326168
rect 311678 326080 311858 326168
rect 311966 326080 312146 326168
rect 312254 326080 312434 326168
rect 312542 326080 312722 326168
rect 312830 326080 313010 326168
rect 325310 326080 325490 326168
rect 325598 326080 325778 326168
rect 325886 326080 326066 326168
rect 326174 326080 326354 326168
rect 326462 326080 326642 326168
rect 326750 326080 326930 326168
rect 327038 326080 327218 326168
rect 327326 326080 327506 326168
rect 339806 326080 339986 326168
rect 340094 326080 340274 326168
rect 340382 326080 340562 326168
rect 340670 326080 340850 326168
rect 340958 326080 341138 326168
rect 341246 326080 341426 326168
rect 341534 326080 341714 326168
rect 341822 326080 342002 326168
rect 354302 326080 354482 326168
rect 354590 326080 354770 326168
rect 354878 326080 355058 326168
rect 355166 326080 355346 326168
rect 355454 326080 355634 326168
rect 355742 326080 355922 326168
rect 356030 326080 356210 326168
rect 356318 326080 356498 326168
rect 368798 326080 368978 326168
rect 369086 326080 369266 326168
rect 369374 326080 369554 326168
rect 369662 326080 369842 326168
rect 369950 326080 370130 326168
rect 370238 326080 370418 326168
rect 370526 326080 370706 326168
rect 370814 326080 370994 326168
rect 383294 326080 383474 326168
rect 383582 326080 383762 326168
rect 383870 326080 384050 326168
rect 384158 326080 384338 326168
rect 384446 326080 384626 326168
rect 384734 326080 384914 326168
rect 385022 326080 385202 326168
rect 385310 326080 385490 326168
rect 397790 326080 397970 326168
rect 398078 326080 398258 326168
rect 398366 326080 398546 326168
rect 398654 326080 398834 326168
rect 398942 326080 399122 326168
rect 399230 326080 399410 326168
rect 399518 326080 399698 326168
rect 399806 326080 399986 326168
rect 412286 326080 412466 326168
rect 412574 326080 412754 326168
rect 412862 326080 413042 326168
rect 413150 326080 413330 326168
rect 413438 326080 413618 326168
rect 413726 326080 413906 326168
rect 414014 326080 414194 326168
rect 414302 326080 414482 326168
rect 426782 326080 426962 326168
rect 427070 326080 427250 326168
rect 427358 326080 427538 326168
rect 427646 326080 427826 326168
rect 427934 326080 428114 326168
rect 428222 326080 428402 326168
rect 428510 326080 428690 326168
rect 428798 326080 428978 326168
rect 441278 326080 441458 326168
rect 441566 326080 441746 326168
rect 441854 326080 442034 326168
rect 442142 326080 442322 326168
rect 442430 326080 442610 326168
rect 442718 326080 442898 326168
rect 443006 326080 443186 326168
rect 443294 326080 443474 326168
rect 455774 326080 455954 326168
rect 456062 326080 456242 326168
rect 456350 326080 456530 326168
rect 456638 326080 456818 326168
rect 456926 326080 457106 326168
rect 457214 326080 457394 326168
rect 457502 326080 457682 326168
rect 457790 326080 457970 326168
rect 180350 311928 180530 312016
rect 180638 311928 180818 312016
rect 180926 311928 181106 312016
rect 181214 311928 181394 312016
rect 181502 311928 181682 312016
rect 181790 311928 181970 312016
rect 182078 311928 182258 312016
rect 182366 311928 182546 312016
rect 194846 311928 195026 312016
rect 195134 311928 195314 312016
rect 195422 311928 195602 312016
rect 195710 311928 195890 312016
rect 195998 311928 196178 312016
rect 196286 311928 196466 312016
rect 196574 311928 196754 312016
rect 196862 311928 197042 312016
rect 209342 311928 209522 312016
rect 209630 311928 209810 312016
rect 209918 311928 210098 312016
rect 210206 311928 210386 312016
rect 210494 311928 210674 312016
rect 210782 311928 210962 312016
rect 211070 311928 211250 312016
rect 211358 311928 211538 312016
rect 223838 311928 224018 312016
rect 224126 311928 224306 312016
rect 224414 311928 224594 312016
rect 224702 311928 224882 312016
rect 224990 311928 225170 312016
rect 225278 311928 225458 312016
rect 225566 311928 225746 312016
rect 225854 311928 226034 312016
rect 238334 311928 238514 312016
rect 238622 311928 238802 312016
rect 238910 311928 239090 312016
rect 239198 311928 239378 312016
rect 239486 311928 239666 312016
rect 239774 311928 239954 312016
rect 240062 311928 240242 312016
rect 240350 311928 240530 312016
rect 252830 311928 253010 312016
rect 253118 311928 253298 312016
rect 253406 311928 253586 312016
rect 253694 311928 253874 312016
rect 253982 311928 254162 312016
rect 254270 311928 254450 312016
rect 254558 311928 254738 312016
rect 254846 311928 255026 312016
rect 267326 311928 267506 312016
rect 267614 311928 267794 312016
rect 267902 311928 268082 312016
rect 268190 311928 268370 312016
rect 268478 311928 268658 312016
rect 268766 311928 268946 312016
rect 269054 311928 269234 312016
rect 269342 311928 269522 312016
rect 281822 311928 282002 312016
rect 282110 311928 282290 312016
rect 282398 311928 282578 312016
rect 282686 311928 282866 312016
rect 282974 311928 283154 312016
rect 283262 311928 283442 312016
rect 283550 311928 283730 312016
rect 283838 311928 284018 312016
rect 296318 311928 296498 312016
rect 296606 311928 296786 312016
rect 296894 311928 297074 312016
rect 297182 311928 297362 312016
rect 297470 311928 297650 312016
rect 297758 311928 297938 312016
rect 298046 311928 298226 312016
rect 298334 311928 298514 312016
rect 310814 311928 310994 312016
rect 311102 311928 311282 312016
rect 311390 311928 311570 312016
rect 311678 311928 311858 312016
rect 311966 311928 312146 312016
rect 312254 311928 312434 312016
rect 312542 311928 312722 312016
rect 312830 311928 313010 312016
rect 325310 311928 325490 312016
rect 325598 311928 325778 312016
rect 325886 311928 326066 312016
rect 326174 311928 326354 312016
rect 326462 311928 326642 312016
rect 326750 311928 326930 312016
rect 327038 311928 327218 312016
rect 327326 311928 327506 312016
rect 339806 311928 339986 312016
rect 340094 311928 340274 312016
rect 340382 311928 340562 312016
rect 340670 311928 340850 312016
rect 340958 311928 341138 312016
rect 341246 311928 341426 312016
rect 341534 311928 341714 312016
rect 341822 311928 342002 312016
rect 354302 311928 354482 312016
rect 354590 311928 354770 312016
rect 354878 311928 355058 312016
rect 355166 311928 355346 312016
rect 355454 311928 355634 312016
rect 355742 311928 355922 312016
rect 356030 311928 356210 312016
rect 356318 311928 356498 312016
rect 368798 311928 368978 312016
rect 369086 311928 369266 312016
rect 369374 311928 369554 312016
rect 369662 311928 369842 312016
rect 369950 311928 370130 312016
rect 370238 311928 370418 312016
rect 370526 311928 370706 312016
rect 370814 311928 370994 312016
rect 383294 311928 383474 312016
rect 383582 311928 383762 312016
rect 383870 311928 384050 312016
rect 384158 311928 384338 312016
rect 384446 311928 384626 312016
rect 384734 311928 384914 312016
rect 385022 311928 385202 312016
rect 385310 311928 385490 312016
rect 397790 311928 397970 312016
rect 398078 311928 398258 312016
rect 398366 311928 398546 312016
rect 398654 311928 398834 312016
rect 398942 311928 399122 312016
rect 399230 311928 399410 312016
rect 399518 311928 399698 312016
rect 399806 311928 399986 312016
rect 412286 311928 412466 312016
rect 412574 311928 412754 312016
rect 412862 311928 413042 312016
rect 413150 311928 413330 312016
rect 413438 311928 413618 312016
rect 413726 311928 413906 312016
rect 414014 311928 414194 312016
rect 414302 311928 414482 312016
rect 426782 311928 426962 312016
rect 427070 311928 427250 312016
rect 427358 311928 427538 312016
rect 427646 311928 427826 312016
rect 427934 311928 428114 312016
rect 428222 311928 428402 312016
rect 428510 311928 428690 312016
rect 428798 311928 428978 312016
rect 441278 311928 441458 312016
rect 441566 311928 441746 312016
rect 441854 311928 442034 312016
rect 442142 311928 442322 312016
rect 442430 311928 442610 312016
rect 442718 311928 442898 312016
rect 443006 311928 443186 312016
rect 443294 311928 443474 312016
rect 455774 311928 455954 312016
rect 456062 311928 456242 312016
rect 456350 311928 456530 312016
rect 456638 311928 456818 312016
rect 456926 311928 457106 312016
rect 457214 311928 457394 312016
rect 457502 311928 457682 312016
rect 457790 311928 457970 312016
rect 180350 311712 180530 311800
rect 180638 311712 180818 311800
rect 180926 311712 181106 311800
rect 181214 311712 181394 311800
rect 181502 311712 181682 311800
rect 181790 311712 181970 311800
rect 182078 311712 182258 311800
rect 182366 311712 182546 311800
rect 194846 311712 195026 311800
rect 195134 311712 195314 311800
rect 195422 311712 195602 311800
rect 195710 311712 195890 311800
rect 195998 311712 196178 311800
rect 196286 311712 196466 311800
rect 196574 311712 196754 311800
rect 196862 311712 197042 311800
rect 209342 311712 209522 311800
rect 209630 311712 209810 311800
rect 209918 311712 210098 311800
rect 210206 311712 210386 311800
rect 210494 311712 210674 311800
rect 210782 311712 210962 311800
rect 211070 311712 211250 311800
rect 211358 311712 211538 311800
rect 223838 311712 224018 311800
rect 224126 311712 224306 311800
rect 224414 311712 224594 311800
rect 224702 311712 224882 311800
rect 224990 311712 225170 311800
rect 225278 311712 225458 311800
rect 225566 311712 225746 311800
rect 225854 311712 226034 311800
rect 238334 311712 238514 311800
rect 238622 311712 238802 311800
rect 238910 311712 239090 311800
rect 239198 311712 239378 311800
rect 239486 311712 239666 311800
rect 239774 311712 239954 311800
rect 240062 311712 240242 311800
rect 240350 311712 240530 311800
rect 252830 311712 253010 311800
rect 253118 311712 253298 311800
rect 253406 311712 253586 311800
rect 253694 311712 253874 311800
rect 253982 311712 254162 311800
rect 254270 311712 254450 311800
rect 254558 311712 254738 311800
rect 254846 311712 255026 311800
rect 267326 311712 267506 311800
rect 267614 311712 267794 311800
rect 267902 311712 268082 311800
rect 268190 311712 268370 311800
rect 268478 311712 268658 311800
rect 268766 311712 268946 311800
rect 269054 311712 269234 311800
rect 269342 311712 269522 311800
rect 281822 311712 282002 311800
rect 282110 311712 282290 311800
rect 282398 311712 282578 311800
rect 282686 311712 282866 311800
rect 282974 311712 283154 311800
rect 283262 311712 283442 311800
rect 283550 311712 283730 311800
rect 283838 311712 284018 311800
rect 296318 311712 296498 311800
rect 296606 311712 296786 311800
rect 296894 311712 297074 311800
rect 297182 311712 297362 311800
rect 297470 311712 297650 311800
rect 297758 311712 297938 311800
rect 298046 311712 298226 311800
rect 298334 311712 298514 311800
rect 310814 311712 310994 311800
rect 311102 311712 311282 311800
rect 311390 311712 311570 311800
rect 311678 311712 311858 311800
rect 311966 311712 312146 311800
rect 312254 311712 312434 311800
rect 312542 311712 312722 311800
rect 312830 311712 313010 311800
rect 325310 311712 325490 311800
rect 325598 311712 325778 311800
rect 325886 311712 326066 311800
rect 326174 311712 326354 311800
rect 326462 311712 326642 311800
rect 326750 311712 326930 311800
rect 327038 311712 327218 311800
rect 327326 311712 327506 311800
rect 339806 311712 339986 311800
rect 340094 311712 340274 311800
rect 340382 311712 340562 311800
rect 340670 311712 340850 311800
rect 340958 311712 341138 311800
rect 341246 311712 341426 311800
rect 341534 311712 341714 311800
rect 341822 311712 342002 311800
rect 354302 311712 354482 311800
rect 354590 311712 354770 311800
rect 354878 311712 355058 311800
rect 355166 311712 355346 311800
rect 355454 311712 355634 311800
rect 355742 311712 355922 311800
rect 356030 311712 356210 311800
rect 356318 311712 356498 311800
rect 368798 311712 368978 311800
rect 369086 311712 369266 311800
rect 369374 311712 369554 311800
rect 369662 311712 369842 311800
rect 369950 311712 370130 311800
rect 370238 311712 370418 311800
rect 370526 311712 370706 311800
rect 370814 311712 370994 311800
rect 383294 311712 383474 311800
rect 383582 311712 383762 311800
rect 383870 311712 384050 311800
rect 384158 311712 384338 311800
rect 384446 311712 384626 311800
rect 384734 311712 384914 311800
rect 385022 311712 385202 311800
rect 385310 311712 385490 311800
rect 397790 311712 397970 311800
rect 398078 311712 398258 311800
rect 398366 311712 398546 311800
rect 398654 311712 398834 311800
rect 398942 311712 399122 311800
rect 399230 311712 399410 311800
rect 399518 311712 399698 311800
rect 399806 311712 399986 311800
rect 412286 311712 412466 311800
rect 412574 311712 412754 311800
rect 412862 311712 413042 311800
rect 413150 311712 413330 311800
rect 413438 311712 413618 311800
rect 413726 311712 413906 311800
rect 414014 311712 414194 311800
rect 414302 311712 414482 311800
rect 426782 311712 426962 311800
rect 427070 311712 427250 311800
rect 427358 311712 427538 311800
rect 427646 311712 427826 311800
rect 427934 311712 428114 311800
rect 428222 311712 428402 311800
rect 428510 311712 428690 311800
rect 428798 311712 428978 311800
rect 441278 311712 441458 311800
rect 441566 311712 441746 311800
rect 441854 311712 442034 311800
rect 442142 311712 442322 311800
rect 442430 311712 442610 311800
rect 442718 311712 442898 311800
rect 443006 311712 443186 311800
rect 443294 311712 443474 311800
rect 455774 311712 455954 311800
rect 456062 311712 456242 311800
rect 456350 311712 456530 311800
rect 456638 311712 456818 311800
rect 456926 311712 457106 311800
rect 457214 311712 457394 311800
rect 457502 311712 457682 311800
rect 457790 311712 457970 311800
rect 180350 311236 180530 311324
rect 180638 311236 180818 311324
rect 180926 311236 181106 311324
rect 181214 311236 181394 311324
rect 181502 311236 181682 311324
rect 181790 311236 181970 311324
rect 182078 311236 182258 311324
rect 182366 311236 182546 311324
rect 194846 311236 195026 311324
rect 195134 311236 195314 311324
rect 195422 311236 195602 311324
rect 195710 311236 195890 311324
rect 195998 311236 196178 311324
rect 196286 311236 196466 311324
rect 196574 311236 196754 311324
rect 196862 311236 197042 311324
rect 209342 311236 209522 311324
rect 209630 311236 209810 311324
rect 209918 311236 210098 311324
rect 210206 311236 210386 311324
rect 210494 311236 210674 311324
rect 210782 311236 210962 311324
rect 211070 311236 211250 311324
rect 211358 311236 211538 311324
rect 223838 311236 224018 311324
rect 224126 311236 224306 311324
rect 224414 311236 224594 311324
rect 224702 311236 224882 311324
rect 224990 311236 225170 311324
rect 225278 311236 225458 311324
rect 225566 311236 225746 311324
rect 225854 311236 226034 311324
rect 238334 311236 238514 311324
rect 238622 311236 238802 311324
rect 238910 311236 239090 311324
rect 239198 311236 239378 311324
rect 239486 311236 239666 311324
rect 239774 311236 239954 311324
rect 240062 311236 240242 311324
rect 240350 311236 240530 311324
rect 252830 311236 253010 311324
rect 253118 311236 253298 311324
rect 253406 311236 253586 311324
rect 253694 311236 253874 311324
rect 253982 311236 254162 311324
rect 254270 311236 254450 311324
rect 254558 311236 254738 311324
rect 254846 311236 255026 311324
rect 267326 311236 267506 311324
rect 267614 311236 267794 311324
rect 267902 311236 268082 311324
rect 268190 311236 268370 311324
rect 268478 311236 268658 311324
rect 268766 311236 268946 311324
rect 269054 311236 269234 311324
rect 269342 311236 269522 311324
rect 281822 311236 282002 311324
rect 282110 311236 282290 311324
rect 282398 311236 282578 311324
rect 282686 311236 282866 311324
rect 282974 311236 283154 311324
rect 283262 311236 283442 311324
rect 283550 311236 283730 311324
rect 283838 311236 284018 311324
rect 296318 311236 296498 311324
rect 296606 311236 296786 311324
rect 296894 311236 297074 311324
rect 297182 311236 297362 311324
rect 297470 311236 297650 311324
rect 297758 311236 297938 311324
rect 298046 311236 298226 311324
rect 298334 311236 298514 311324
rect 310814 311236 310994 311324
rect 311102 311236 311282 311324
rect 311390 311236 311570 311324
rect 311678 311236 311858 311324
rect 311966 311236 312146 311324
rect 312254 311236 312434 311324
rect 312542 311236 312722 311324
rect 312830 311236 313010 311324
rect 325310 311236 325490 311324
rect 325598 311236 325778 311324
rect 325886 311236 326066 311324
rect 326174 311236 326354 311324
rect 326462 311236 326642 311324
rect 326750 311236 326930 311324
rect 327038 311236 327218 311324
rect 327326 311236 327506 311324
rect 339806 311236 339986 311324
rect 340094 311236 340274 311324
rect 340382 311236 340562 311324
rect 340670 311236 340850 311324
rect 340958 311236 341138 311324
rect 341246 311236 341426 311324
rect 341534 311236 341714 311324
rect 341822 311236 342002 311324
rect 354302 311236 354482 311324
rect 354590 311236 354770 311324
rect 354878 311236 355058 311324
rect 355166 311236 355346 311324
rect 355454 311236 355634 311324
rect 355742 311236 355922 311324
rect 356030 311236 356210 311324
rect 356318 311236 356498 311324
rect 368798 311236 368978 311324
rect 369086 311236 369266 311324
rect 369374 311236 369554 311324
rect 369662 311236 369842 311324
rect 369950 311236 370130 311324
rect 370238 311236 370418 311324
rect 370526 311236 370706 311324
rect 370814 311236 370994 311324
rect 383294 311236 383474 311324
rect 383582 311236 383762 311324
rect 383870 311236 384050 311324
rect 384158 311236 384338 311324
rect 384446 311236 384626 311324
rect 384734 311236 384914 311324
rect 385022 311236 385202 311324
rect 385310 311236 385490 311324
rect 397790 311236 397970 311324
rect 398078 311236 398258 311324
rect 398366 311236 398546 311324
rect 398654 311236 398834 311324
rect 398942 311236 399122 311324
rect 399230 311236 399410 311324
rect 399518 311236 399698 311324
rect 399806 311236 399986 311324
rect 412286 311236 412466 311324
rect 412574 311236 412754 311324
rect 412862 311236 413042 311324
rect 413150 311236 413330 311324
rect 413438 311236 413618 311324
rect 413726 311236 413906 311324
rect 414014 311236 414194 311324
rect 414302 311236 414482 311324
rect 426782 311236 426962 311324
rect 427070 311236 427250 311324
rect 427358 311236 427538 311324
rect 427646 311236 427826 311324
rect 427934 311236 428114 311324
rect 428222 311236 428402 311324
rect 428510 311236 428690 311324
rect 428798 311236 428978 311324
rect 441278 311236 441458 311324
rect 441566 311236 441746 311324
rect 441854 311236 442034 311324
rect 442142 311236 442322 311324
rect 442430 311236 442610 311324
rect 442718 311236 442898 311324
rect 443006 311236 443186 311324
rect 443294 311236 443474 311324
rect 455774 311236 455954 311324
rect 456062 311236 456242 311324
rect 456350 311236 456530 311324
rect 456638 311236 456818 311324
rect 456926 311236 457106 311324
rect 457214 311236 457394 311324
rect 457502 311236 457682 311324
rect 457790 311236 457970 311324
rect 180350 311020 180530 311108
rect 180638 311020 180818 311108
rect 180926 311020 181106 311108
rect 181214 311020 181394 311108
rect 181502 311020 181682 311108
rect 181790 311020 181970 311108
rect 182078 311020 182258 311108
rect 182366 311020 182546 311108
rect 194846 311020 195026 311108
rect 195134 311020 195314 311108
rect 195422 311020 195602 311108
rect 195710 311020 195890 311108
rect 195998 311020 196178 311108
rect 196286 311020 196466 311108
rect 196574 311020 196754 311108
rect 196862 311020 197042 311108
rect 209342 311020 209522 311108
rect 209630 311020 209810 311108
rect 209918 311020 210098 311108
rect 210206 311020 210386 311108
rect 210494 311020 210674 311108
rect 210782 311020 210962 311108
rect 211070 311020 211250 311108
rect 211358 311020 211538 311108
rect 223838 311020 224018 311108
rect 224126 311020 224306 311108
rect 224414 311020 224594 311108
rect 224702 311020 224882 311108
rect 224990 311020 225170 311108
rect 225278 311020 225458 311108
rect 225566 311020 225746 311108
rect 225854 311020 226034 311108
rect 238334 311020 238514 311108
rect 238622 311020 238802 311108
rect 238910 311020 239090 311108
rect 239198 311020 239378 311108
rect 239486 311020 239666 311108
rect 239774 311020 239954 311108
rect 240062 311020 240242 311108
rect 240350 311020 240530 311108
rect 252830 311020 253010 311108
rect 253118 311020 253298 311108
rect 253406 311020 253586 311108
rect 253694 311020 253874 311108
rect 253982 311020 254162 311108
rect 254270 311020 254450 311108
rect 254558 311020 254738 311108
rect 254846 311020 255026 311108
rect 267326 311020 267506 311108
rect 267614 311020 267794 311108
rect 267902 311020 268082 311108
rect 268190 311020 268370 311108
rect 268478 311020 268658 311108
rect 268766 311020 268946 311108
rect 269054 311020 269234 311108
rect 269342 311020 269522 311108
rect 281822 311020 282002 311108
rect 282110 311020 282290 311108
rect 282398 311020 282578 311108
rect 282686 311020 282866 311108
rect 282974 311020 283154 311108
rect 283262 311020 283442 311108
rect 283550 311020 283730 311108
rect 283838 311020 284018 311108
rect 296318 311020 296498 311108
rect 296606 311020 296786 311108
rect 296894 311020 297074 311108
rect 297182 311020 297362 311108
rect 297470 311020 297650 311108
rect 297758 311020 297938 311108
rect 298046 311020 298226 311108
rect 298334 311020 298514 311108
rect 310814 311020 310994 311108
rect 311102 311020 311282 311108
rect 311390 311020 311570 311108
rect 311678 311020 311858 311108
rect 311966 311020 312146 311108
rect 312254 311020 312434 311108
rect 312542 311020 312722 311108
rect 312830 311020 313010 311108
rect 325310 311020 325490 311108
rect 325598 311020 325778 311108
rect 325886 311020 326066 311108
rect 326174 311020 326354 311108
rect 326462 311020 326642 311108
rect 326750 311020 326930 311108
rect 327038 311020 327218 311108
rect 327326 311020 327506 311108
rect 339806 311020 339986 311108
rect 340094 311020 340274 311108
rect 340382 311020 340562 311108
rect 340670 311020 340850 311108
rect 340958 311020 341138 311108
rect 341246 311020 341426 311108
rect 341534 311020 341714 311108
rect 341822 311020 342002 311108
rect 354302 311020 354482 311108
rect 354590 311020 354770 311108
rect 354878 311020 355058 311108
rect 355166 311020 355346 311108
rect 355454 311020 355634 311108
rect 355742 311020 355922 311108
rect 356030 311020 356210 311108
rect 356318 311020 356498 311108
rect 368798 311020 368978 311108
rect 369086 311020 369266 311108
rect 369374 311020 369554 311108
rect 369662 311020 369842 311108
rect 369950 311020 370130 311108
rect 370238 311020 370418 311108
rect 370526 311020 370706 311108
rect 370814 311020 370994 311108
rect 383294 311020 383474 311108
rect 383582 311020 383762 311108
rect 383870 311020 384050 311108
rect 384158 311020 384338 311108
rect 384446 311020 384626 311108
rect 384734 311020 384914 311108
rect 385022 311020 385202 311108
rect 385310 311020 385490 311108
rect 397790 311020 397970 311108
rect 398078 311020 398258 311108
rect 398366 311020 398546 311108
rect 398654 311020 398834 311108
rect 398942 311020 399122 311108
rect 399230 311020 399410 311108
rect 399518 311020 399698 311108
rect 399806 311020 399986 311108
rect 412286 311020 412466 311108
rect 412574 311020 412754 311108
rect 412862 311020 413042 311108
rect 413150 311020 413330 311108
rect 413438 311020 413618 311108
rect 413726 311020 413906 311108
rect 414014 311020 414194 311108
rect 414302 311020 414482 311108
rect 426782 311020 426962 311108
rect 427070 311020 427250 311108
rect 427358 311020 427538 311108
rect 427646 311020 427826 311108
rect 427934 311020 428114 311108
rect 428222 311020 428402 311108
rect 428510 311020 428690 311108
rect 428798 311020 428978 311108
rect 441278 311020 441458 311108
rect 441566 311020 441746 311108
rect 441854 311020 442034 311108
rect 442142 311020 442322 311108
rect 442430 311020 442610 311108
rect 442718 311020 442898 311108
rect 443006 311020 443186 311108
rect 443294 311020 443474 311108
rect 455774 311020 455954 311108
rect 456062 311020 456242 311108
rect 456350 311020 456530 311108
rect 456638 311020 456818 311108
rect 456926 311020 457106 311108
rect 457214 311020 457394 311108
rect 457502 311020 457682 311108
rect 457790 311020 457970 311108
rect 180350 296868 180530 296956
rect 180638 296868 180818 296956
rect 180926 296868 181106 296956
rect 181214 296868 181394 296956
rect 181502 296868 181682 296956
rect 181790 296868 181970 296956
rect 182078 296868 182258 296956
rect 182366 296868 182546 296956
rect 194846 296868 195026 296956
rect 195134 296868 195314 296956
rect 195422 296868 195602 296956
rect 195710 296868 195890 296956
rect 195998 296868 196178 296956
rect 196286 296868 196466 296956
rect 196574 296868 196754 296956
rect 196862 296868 197042 296956
rect 209342 296868 209522 296956
rect 209630 296868 209810 296956
rect 209918 296868 210098 296956
rect 210206 296868 210386 296956
rect 210494 296868 210674 296956
rect 210782 296868 210962 296956
rect 211070 296868 211250 296956
rect 211358 296868 211538 296956
rect 223838 296868 224018 296956
rect 224126 296868 224306 296956
rect 224414 296868 224594 296956
rect 224702 296868 224882 296956
rect 224990 296868 225170 296956
rect 225278 296868 225458 296956
rect 225566 296868 225746 296956
rect 225854 296868 226034 296956
rect 238334 296868 238514 296956
rect 238622 296868 238802 296956
rect 238910 296868 239090 296956
rect 239198 296868 239378 296956
rect 239486 296868 239666 296956
rect 239774 296868 239954 296956
rect 240062 296868 240242 296956
rect 240350 296868 240530 296956
rect 252830 296868 253010 296956
rect 253118 296868 253298 296956
rect 253406 296868 253586 296956
rect 253694 296868 253874 296956
rect 253982 296868 254162 296956
rect 254270 296868 254450 296956
rect 254558 296868 254738 296956
rect 254846 296868 255026 296956
rect 267326 296868 267506 296956
rect 267614 296868 267794 296956
rect 267902 296868 268082 296956
rect 268190 296868 268370 296956
rect 268478 296868 268658 296956
rect 268766 296868 268946 296956
rect 269054 296868 269234 296956
rect 269342 296868 269522 296956
rect 281822 296868 282002 296956
rect 282110 296868 282290 296956
rect 282398 296868 282578 296956
rect 282686 296868 282866 296956
rect 282974 296868 283154 296956
rect 283262 296868 283442 296956
rect 283550 296868 283730 296956
rect 283838 296868 284018 296956
rect 296318 296868 296498 296956
rect 296606 296868 296786 296956
rect 296894 296868 297074 296956
rect 297182 296868 297362 296956
rect 297470 296868 297650 296956
rect 297758 296868 297938 296956
rect 298046 296868 298226 296956
rect 298334 296868 298514 296956
rect 310814 296868 310994 296956
rect 311102 296868 311282 296956
rect 311390 296868 311570 296956
rect 311678 296868 311858 296956
rect 311966 296868 312146 296956
rect 312254 296868 312434 296956
rect 312542 296868 312722 296956
rect 312830 296868 313010 296956
rect 325310 296868 325490 296956
rect 325598 296868 325778 296956
rect 325886 296868 326066 296956
rect 326174 296868 326354 296956
rect 326462 296868 326642 296956
rect 326750 296868 326930 296956
rect 327038 296868 327218 296956
rect 327326 296868 327506 296956
rect 339806 296868 339986 296956
rect 340094 296868 340274 296956
rect 340382 296868 340562 296956
rect 340670 296868 340850 296956
rect 340958 296868 341138 296956
rect 341246 296868 341426 296956
rect 341534 296868 341714 296956
rect 341822 296868 342002 296956
rect 354302 296868 354482 296956
rect 354590 296868 354770 296956
rect 354878 296868 355058 296956
rect 355166 296868 355346 296956
rect 355454 296868 355634 296956
rect 355742 296868 355922 296956
rect 356030 296868 356210 296956
rect 356318 296868 356498 296956
rect 368798 296868 368978 296956
rect 369086 296868 369266 296956
rect 369374 296868 369554 296956
rect 369662 296868 369842 296956
rect 369950 296868 370130 296956
rect 370238 296868 370418 296956
rect 370526 296868 370706 296956
rect 370814 296868 370994 296956
rect 383294 296868 383474 296956
rect 383582 296868 383762 296956
rect 383870 296868 384050 296956
rect 384158 296868 384338 296956
rect 384446 296868 384626 296956
rect 384734 296868 384914 296956
rect 385022 296868 385202 296956
rect 385310 296868 385490 296956
rect 397790 296868 397970 296956
rect 398078 296868 398258 296956
rect 398366 296868 398546 296956
rect 398654 296868 398834 296956
rect 398942 296868 399122 296956
rect 399230 296868 399410 296956
rect 399518 296868 399698 296956
rect 399806 296868 399986 296956
rect 412286 296868 412466 296956
rect 412574 296868 412754 296956
rect 412862 296868 413042 296956
rect 413150 296868 413330 296956
rect 413438 296868 413618 296956
rect 413726 296868 413906 296956
rect 414014 296868 414194 296956
rect 414302 296868 414482 296956
rect 426782 296868 426962 296956
rect 427070 296868 427250 296956
rect 427358 296868 427538 296956
rect 427646 296868 427826 296956
rect 427934 296868 428114 296956
rect 428222 296868 428402 296956
rect 428510 296868 428690 296956
rect 428798 296868 428978 296956
rect 441278 296868 441458 296956
rect 441566 296868 441746 296956
rect 441854 296868 442034 296956
rect 442142 296868 442322 296956
rect 442430 296868 442610 296956
rect 442718 296868 442898 296956
rect 443006 296868 443186 296956
rect 443294 296868 443474 296956
rect 455774 296868 455954 296956
rect 456062 296868 456242 296956
rect 456350 296868 456530 296956
rect 456638 296868 456818 296956
rect 456926 296868 457106 296956
rect 457214 296868 457394 296956
rect 457502 296868 457682 296956
rect 457790 296868 457970 296956
rect 180350 296652 180530 296740
rect 180638 296652 180818 296740
rect 180926 296652 181106 296740
rect 181214 296652 181394 296740
rect 181502 296652 181682 296740
rect 181790 296652 181970 296740
rect 182078 296652 182258 296740
rect 182366 296652 182546 296740
rect 194846 296652 195026 296740
rect 195134 296652 195314 296740
rect 195422 296652 195602 296740
rect 195710 296652 195890 296740
rect 195998 296652 196178 296740
rect 196286 296652 196466 296740
rect 196574 296652 196754 296740
rect 196862 296652 197042 296740
rect 209342 296652 209522 296740
rect 209630 296652 209810 296740
rect 209918 296652 210098 296740
rect 210206 296652 210386 296740
rect 210494 296652 210674 296740
rect 210782 296652 210962 296740
rect 211070 296652 211250 296740
rect 211358 296652 211538 296740
rect 223838 296652 224018 296740
rect 224126 296652 224306 296740
rect 224414 296652 224594 296740
rect 224702 296652 224882 296740
rect 224990 296652 225170 296740
rect 225278 296652 225458 296740
rect 225566 296652 225746 296740
rect 225854 296652 226034 296740
rect 238334 296652 238514 296740
rect 238622 296652 238802 296740
rect 238910 296652 239090 296740
rect 239198 296652 239378 296740
rect 239486 296652 239666 296740
rect 239774 296652 239954 296740
rect 240062 296652 240242 296740
rect 240350 296652 240530 296740
rect 252830 296652 253010 296740
rect 253118 296652 253298 296740
rect 253406 296652 253586 296740
rect 253694 296652 253874 296740
rect 253982 296652 254162 296740
rect 254270 296652 254450 296740
rect 254558 296652 254738 296740
rect 254846 296652 255026 296740
rect 267326 296652 267506 296740
rect 267614 296652 267794 296740
rect 267902 296652 268082 296740
rect 268190 296652 268370 296740
rect 268478 296652 268658 296740
rect 268766 296652 268946 296740
rect 269054 296652 269234 296740
rect 269342 296652 269522 296740
rect 281822 296652 282002 296740
rect 282110 296652 282290 296740
rect 282398 296652 282578 296740
rect 282686 296652 282866 296740
rect 282974 296652 283154 296740
rect 283262 296652 283442 296740
rect 283550 296652 283730 296740
rect 283838 296652 284018 296740
rect 296318 296652 296498 296740
rect 296606 296652 296786 296740
rect 296894 296652 297074 296740
rect 297182 296652 297362 296740
rect 297470 296652 297650 296740
rect 297758 296652 297938 296740
rect 298046 296652 298226 296740
rect 298334 296652 298514 296740
rect 310814 296652 310994 296740
rect 311102 296652 311282 296740
rect 311390 296652 311570 296740
rect 311678 296652 311858 296740
rect 311966 296652 312146 296740
rect 312254 296652 312434 296740
rect 312542 296652 312722 296740
rect 312830 296652 313010 296740
rect 325310 296652 325490 296740
rect 325598 296652 325778 296740
rect 325886 296652 326066 296740
rect 326174 296652 326354 296740
rect 326462 296652 326642 296740
rect 326750 296652 326930 296740
rect 327038 296652 327218 296740
rect 327326 296652 327506 296740
rect 339806 296652 339986 296740
rect 340094 296652 340274 296740
rect 340382 296652 340562 296740
rect 340670 296652 340850 296740
rect 340958 296652 341138 296740
rect 341246 296652 341426 296740
rect 341534 296652 341714 296740
rect 341822 296652 342002 296740
rect 354302 296652 354482 296740
rect 354590 296652 354770 296740
rect 354878 296652 355058 296740
rect 355166 296652 355346 296740
rect 355454 296652 355634 296740
rect 355742 296652 355922 296740
rect 356030 296652 356210 296740
rect 356318 296652 356498 296740
rect 368798 296652 368978 296740
rect 369086 296652 369266 296740
rect 369374 296652 369554 296740
rect 369662 296652 369842 296740
rect 369950 296652 370130 296740
rect 370238 296652 370418 296740
rect 370526 296652 370706 296740
rect 370814 296652 370994 296740
rect 383294 296652 383474 296740
rect 383582 296652 383762 296740
rect 383870 296652 384050 296740
rect 384158 296652 384338 296740
rect 384446 296652 384626 296740
rect 384734 296652 384914 296740
rect 385022 296652 385202 296740
rect 385310 296652 385490 296740
rect 397790 296652 397970 296740
rect 398078 296652 398258 296740
rect 398366 296652 398546 296740
rect 398654 296652 398834 296740
rect 398942 296652 399122 296740
rect 399230 296652 399410 296740
rect 399518 296652 399698 296740
rect 399806 296652 399986 296740
rect 412286 296652 412466 296740
rect 412574 296652 412754 296740
rect 412862 296652 413042 296740
rect 413150 296652 413330 296740
rect 413438 296652 413618 296740
rect 413726 296652 413906 296740
rect 414014 296652 414194 296740
rect 414302 296652 414482 296740
rect 426782 296652 426962 296740
rect 427070 296652 427250 296740
rect 427358 296652 427538 296740
rect 427646 296652 427826 296740
rect 427934 296652 428114 296740
rect 428222 296652 428402 296740
rect 428510 296652 428690 296740
rect 428798 296652 428978 296740
rect 441278 296652 441458 296740
rect 441566 296652 441746 296740
rect 441854 296652 442034 296740
rect 442142 296652 442322 296740
rect 442430 296652 442610 296740
rect 442718 296652 442898 296740
rect 443006 296652 443186 296740
rect 443294 296652 443474 296740
rect 455774 296652 455954 296740
rect 456062 296652 456242 296740
rect 456350 296652 456530 296740
rect 456638 296652 456818 296740
rect 456926 296652 457106 296740
rect 457214 296652 457394 296740
rect 457502 296652 457682 296740
rect 457790 296652 457970 296740
rect 180350 296176 180530 296264
rect 180638 296176 180818 296264
rect 180926 296176 181106 296264
rect 181214 296176 181394 296264
rect 181502 296176 181682 296264
rect 181790 296176 181970 296264
rect 182078 296176 182258 296264
rect 182366 296176 182546 296264
rect 194846 296176 195026 296264
rect 195134 296176 195314 296264
rect 195422 296176 195602 296264
rect 195710 296176 195890 296264
rect 195998 296176 196178 296264
rect 196286 296176 196466 296264
rect 196574 296176 196754 296264
rect 196862 296176 197042 296264
rect 209342 296176 209522 296264
rect 209630 296176 209810 296264
rect 209918 296176 210098 296264
rect 210206 296176 210386 296264
rect 210494 296176 210674 296264
rect 210782 296176 210962 296264
rect 211070 296176 211250 296264
rect 211358 296176 211538 296264
rect 223838 296176 224018 296264
rect 224126 296176 224306 296264
rect 224414 296176 224594 296264
rect 224702 296176 224882 296264
rect 224990 296176 225170 296264
rect 225278 296176 225458 296264
rect 225566 296176 225746 296264
rect 225854 296176 226034 296264
rect 238334 296176 238514 296264
rect 238622 296176 238802 296264
rect 238910 296176 239090 296264
rect 239198 296176 239378 296264
rect 239486 296176 239666 296264
rect 239774 296176 239954 296264
rect 240062 296176 240242 296264
rect 240350 296176 240530 296264
rect 252830 296176 253010 296264
rect 253118 296176 253298 296264
rect 253406 296176 253586 296264
rect 253694 296176 253874 296264
rect 253982 296176 254162 296264
rect 254270 296176 254450 296264
rect 254558 296176 254738 296264
rect 254846 296176 255026 296264
rect 267326 296176 267506 296264
rect 267614 296176 267794 296264
rect 267902 296176 268082 296264
rect 268190 296176 268370 296264
rect 268478 296176 268658 296264
rect 268766 296176 268946 296264
rect 269054 296176 269234 296264
rect 269342 296176 269522 296264
rect 281822 296176 282002 296264
rect 282110 296176 282290 296264
rect 282398 296176 282578 296264
rect 282686 296176 282866 296264
rect 282974 296176 283154 296264
rect 283262 296176 283442 296264
rect 283550 296176 283730 296264
rect 283838 296176 284018 296264
rect 296318 296176 296498 296264
rect 296606 296176 296786 296264
rect 296894 296176 297074 296264
rect 297182 296176 297362 296264
rect 297470 296176 297650 296264
rect 297758 296176 297938 296264
rect 298046 296176 298226 296264
rect 298334 296176 298514 296264
rect 310814 296176 310994 296264
rect 311102 296176 311282 296264
rect 311390 296176 311570 296264
rect 311678 296176 311858 296264
rect 311966 296176 312146 296264
rect 312254 296176 312434 296264
rect 312542 296176 312722 296264
rect 312830 296176 313010 296264
rect 325310 296176 325490 296264
rect 325598 296176 325778 296264
rect 325886 296176 326066 296264
rect 326174 296176 326354 296264
rect 326462 296176 326642 296264
rect 326750 296176 326930 296264
rect 327038 296176 327218 296264
rect 327326 296176 327506 296264
rect 339806 296176 339986 296264
rect 340094 296176 340274 296264
rect 340382 296176 340562 296264
rect 340670 296176 340850 296264
rect 340958 296176 341138 296264
rect 341246 296176 341426 296264
rect 341534 296176 341714 296264
rect 341822 296176 342002 296264
rect 354302 296176 354482 296264
rect 354590 296176 354770 296264
rect 354878 296176 355058 296264
rect 355166 296176 355346 296264
rect 355454 296176 355634 296264
rect 355742 296176 355922 296264
rect 356030 296176 356210 296264
rect 356318 296176 356498 296264
rect 368798 296176 368978 296264
rect 369086 296176 369266 296264
rect 369374 296176 369554 296264
rect 369662 296176 369842 296264
rect 369950 296176 370130 296264
rect 370238 296176 370418 296264
rect 370526 296176 370706 296264
rect 370814 296176 370994 296264
rect 383294 296176 383474 296264
rect 383582 296176 383762 296264
rect 383870 296176 384050 296264
rect 384158 296176 384338 296264
rect 384446 296176 384626 296264
rect 384734 296176 384914 296264
rect 385022 296176 385202 296264
rect 385310 296176 385490 296264
rect 397790 296176 397970 296264
rect 398078 296176 398258 296264
rect 398366 296176 398546 296264
rect 398654 296176 398834 296264
rect 398942 296176 399122 296264
rect 399230 296176 399410 296264
rect 399518 296176 399698 296264
rect 399806 296176 399986 296264
rect 412286 296176 412466 296264
rect 412574 296176 412754 296264
rect 412862 296176 413042 296264
rect 413150 296176 413330 296264
rect 413438 296176 413618 296264
rect 413726 296176 413906 296264
rect 414014 296176 414194 296264
rect 414302 296176 414482 296264
rect 426782 296176 426962 296264
rect 427070 296176 427250 296264
rect 427358 296176 427538 296264
rect 427646 296176 427826 296264
rect 427934 296176 428114 296264
rect 428222 296176 428402 296264
rect 428510 296176 428690 296264
rect 428798 296176 428978 296264
rect 441278 296176 441458 296264
rect 441566 296176 441746 296264
rect 441854 296176 442034 296264
rect 442142 296176 442322 296264
rect 442430 296176 442610 296264
rect 442718 296176 442898 296264
rect 443006 296176 443186 296264
rect 443294 296176 443474 296264
rect 455774 296176 455954 296264
rect 456062 296176 456242 296264
rect 456350 296176 456530 296264
rect 456638 296176 456818 296264
rect 456926 296176 457106 296264
rect 457214 296176 457394 296264
rect 457502 296176 457682 296264
rect 457790 296176 457970 296264
rect 180350 295960 180530 296048
rect 180638 295960 180818 296048
rect 180926 295960 181106 296048
rect 181214 295960 181394 296048
rect 181502 295960 181682 296048
rect 181790 295960 181970 296048
rect 182078 295960 182258 296048
rect 182366 295960 182546 296048
rect 194846 295960 195026 296048
rect 195134 295960 195314 296048
rect 195422 295960 195602 296048
rect 195710 295960 195890 296048
rect 195998 295960 196178 296048
rect 196286 295960 196466 296048
rect 196574 295960 196754 296048
rect 196862 295960 197042 296048
rect 209342 295960 209522 296048
rect 209630 295960 209810 296048
rect 209918 295960 210098 296048
rect 210206 295960 210386 296048
rect 210494 295960 210674 296048
rect 210782 295960 210962 296048
rect 211070 295960 211250 296048
rect 211358 295960 211538 296048
rect 223838 295960 224018 296048
rect 224126 295960 224306 296048
rect 224414 295960 224594 296048
rect 224702 295960 224882 296048
rect 224990 295960 225170 296048
rect 225278 295960 225458 296048
rect 225566 295960 225746 296048
rect 225854 295960 226034 296048
rect 238334 295960 238514 296048
rect 238622 295960 238802 296048
rect 238910 295960 239090 296048
rect 239198 295960 239378 296048
rect 239486 295960 239666 296048
rect 239774 295960 239954 296048
rect 240062 295960 240242 296048
rect 240350 295960 240530 296048
rect 252830 295960 253010 296048
rect 253118 295960 253298 296048
rect 253406 295960 253586 296048
rect 253694 295960 253874 296048
rect 253982 295960 254162 296048
rect 254270 295960 254450 296048
rect 254558 295960 254738 296048
rect 254846 295960 255026 296048
rect 267326 295960 267506 296048
rect 267614 295960 267794 296048
rect 267902 295960 268082 296048
rect 268190 295960 268370 296048
rect 268478 295960 268658 296048
rect 268766 295960 268946 296048
rect 269054 295960 269234 296048
rect 269342 295960 269522 296048
rect 281822 295960 282002 296048
rect 282110 295960 282290 296048
rect 282398 295960 282578 296048
rect 282686 295960 282866 296048
rect 282974 295960 283154 296048
rect 283262 295960 283442 296048
rect 283550 295960 283730 296048
rect 283838 295960 284018 296048
rect 296318 295960 296498 296048
rect 296606 295960 296786 296048
rect 296894 295960 297074 296048
rect 297182 295960 297362 296048
rect 297470 295960 297650 296048
rect 297758 295960 297938 296048
rect 298046 295960 298226 296048
rect 298334 295960 298514 296048
rect 310814 295960 310994 296048
rect 311102 295960 311282 296048
rect 311390 295960 311570 296048
rect 311678 295960 311858 296048
rect 311966 295960 312146 296048
rect 312254 295960 312434 296048
rect 312542 295960 312722 296048
rect 312830 295960 313010 296048
rect 325310 295960 325490 296048
rect 325598 295960 325778 296048
rect 325886 295960 326066 296048
rect 326174 295960 326354 296048
rect 326462 295960 326642 296048
rect 326750 295960 326930 296048
rect 327038 295960 327218 296048
rect 327326 295960 327506 296048
rect 339806 295960 339986 296048
rect 340094 295960 340274 296048
rect 340382 295960 340562 296048
rect 340670 295960 340850 296048
rect 340958 295960 341138 296048
rect 341246 295960 341426 296048
rect 341534 295960 341714 296048
rect 341822 295960 342002 296048
rect 354302 295960 354482 296048
rect 354590 295960 354770 296048
rect 354878 295960 355058 296048
rect 355166 295960 355346 296048
rect 355454 295960 355634 296048
rect 355742 295960 355922 296048
rect 356030 295960 356210 296048
rect 356318 295960 356498 296048
rect 368798 295960 368978 296048
rect 369086 295960 369266 296048
rect 369374 295960 369554 296048
rect 369662 295960 369842 296048
rect 369950 295960 370130 296048
rect 370238 295960 370418 296048
rect 370526 295960 370706 296048
rect 370814 295960 370994 296048
rect 383294 295960 383474 296048
rect 383582 295960 383762 296048
rect 383870 295960 384050 296048
rect 384158 295960 384338 296048
rect 384446 295960 384626 296048
rect 384734 295960 384914 296048
rect 385022 295960 385202 296048
rect 385310 295960 385490 296048
rect 397790 295960 397970 296048
rect 398078 295960 398258 296048
rect 398366 295960 398546 296048
rect 398654 295960 398834 296048
rect 398942 295960 399122 296048
rect 399230 295960 399410 296048
rect 399518 295960 399698 296048
rect 399806 295960 399986 296048
rect 412286 295960 412466 296048
rect 412574 295960 412754 296048
rect 412862 295960 413042 296048
rect 413150 295960 413330 296048
rect 413438 295960 413618 296048
rect 413726 295960 413906 296048
rect 414014 295960 414194 296048
rect 414302 295960 414482 296048
rect 426782 295960 426962 296048
rect 427070 295960 427250 296048
rect 427358 295960 427538 296048
rect 427646 295960 427826 296048
rect 427934 295960 428114 296048
rect 428222 295960 428402 296048
rect 428510 295960 428690 296048
rect 428798 295960 428978 296048
rect 441278 295960 441458 296048
rect 441566 295960 441746 296048
rect 441854 295960 442034 296048
rect 442142 295960 442322 296048
rect 442430 295960 442610 296048
rect 442718 295960 442898 296048
rect 443006 295960 443186 296048
rect 443294 295960 443474 296048
rect 455774 295960 455954 296048
rect 456062 295960 456242 296048
rect 456350 295960 456530 296048
rect 456638 295960 456818 296048
rect 456926 295960 457106 296048
rect 457214 295960 457394 296048
rect 457502 295960 457682 296048
rect 457790 295960 457970 296048
rect 180350 281808 180530 281896
rect 180638 281808 180818 281896
rect 180926 281808 181106 281896
rect 181214 281808 181394 281896
rect 181502 281808 181682 281896
rect 181790 281808 181970 281896
rect 182078 281808 182258 281896
rect 182366 281808 182546 281896
rect 194846 281808 195026 281896
rect 195134 281808 195314 281896
rect 195422 281808 195602 281896
rect 195710 281808 195890 281896
rect 195998 281808 196178 281896
rect 196286 281808 196466 281896
rect 196574 281808 196754 281896
rect 196862 281808 197042 281896
rect 209342 281808 209522 281896
rect 209630 281808 209810 281896
rect 209918 281808 210098 281896
rect 210206 281808 210386 281896
rect 210494 281808 210674 281896
rect 210782 281808 210962 281896
rect 211070 281808 211250 281896
rect 211358 281808 211538 281896
rect 223838 281808 224018 281896
rect 224126 281808 224306 281896
rect 224414 281808 224594 281896
rect 224702 281808 224882 281896
rect 224990 281808 225170 281896
rect 225278 281808 225458 281896
rect 225566 281808 225746 281896
rect 225854 281808 226034 281896
rect 238334 281808 238514 281896
rect 238622 281808 238802 281896
rect 238910 281808 239090 281896
rect 239198 281808 239378 281896
rect 239486 281808 239666 281896
rect 239774 281808 239954 281896
rect 240062 281808 240242 281896
rect 240350 281808 240530 281896
rect 252830 281808 253010 281896
rect 253118 281808 253298 281896
rect 253406 281808 253586 281896
rect 253694 281808 253874 281896
rect 253982 281808 254162 281896
rect 254270 281808 254450 281896
rect 254558 281808 254738 281896
rect 254846 281808 255026 281896
rect 267326 281808 267506 281896
rect 267614 281808 267794 281896
rect 267902 281808 268082 281896
rect 268190 281808 268370 281896
rect 268478 281808 268658 281896
rect 268766 281808 268946 281896
rect 269054 281808 269234 281896
rect 269342 281808 269522 281896
rect 281822 281808 282002 281896
rect 282110 281808 282290 281896
rect 282398 281808 282578 281896
rect 282686 281808 282866 281896
rect 282974 281808 283154 281896
rect 283262 281808 283442 281896
rect 283550 281808 283730 281896
rect 283838 281808 284018 281896
rect 296318 281808 296498 281896
rect 296606 281808 296786 281896
rect 296894 281808 297074 281896
rect 297182 281808 297362 281896
rect 297470 281808 297650 281896
rect 297758 281808 297938 281896
rect 298046 281808 298226 281896
rect 298334 281808 298514 281896
rect 310814 281808 310994 281896
rect 311102 281808 311282 281896
rect 311390 281808 311570 281896
rect 311678 281808 311858 281896
rect 311966 281808 312146 281896
rect 312254 281808 312434 281896
rect 312542 281808 312722 281896
rect 312830 281808 313010 281896
rect 325310 281808 325490 281896
rect 325598 281808 325778 281896
rect 325886 281808 326066 281896
rect 326174 281808 326354 281896
rect 326462 281808 326642 281896
rect 326750 281808 326930 281896
rect 327038 281808 327218 281896
rect 327326 281808 327506 281896
rect 339806 281808 339986 281896
rect 340094 281808 340274 281896
rect 340382 281808 340562 281896
rect 340670 281808 340850 281896
rect 340958 281808 341138 281896
rect 341246 281808 341426 281896
rect 341534 281808 341714 281896
rect 341822 281808 342002 281896
rect 354302 281808 354482 281896
rect 354590 281808 354770 281896
rect 354878 281808 355058 281896
rect 355166 281808 355346 281896
rect 355454 281808 355634 281896
rect 355742 281808 355922 281896
rect 356030 281808 356210 281896
rect 356318 281808 356498 281896
rect 368798 281808 368978 281896
rect 369086 281808 369266 281896
rect 369374 281808 369554 281896
rect 369662 281808 369842 281896
rect 369950 281808 370130 281896
rect 370238 281808 370418 281896
rect 370526 281808 370706 281896
rect 370814 281808 370994 281896
rect 383294 281808 383474 281896
rect 383582 281808 383762 281896
rect 383870 281808 384050 281896
rect 384158 281808 384338 281896
rect 384446 281808 384626 281896
rect 384734 281808 384914 281896
rect 385022 281808 385202 281896
rect 385310 281808 385490 281896
rect 397790 281808 397970 281896
rect 398078 281808 398258 281896
rect 398366 281808 398546 281896
rect 398654 281808 398834 281896
rect 398942 281808 399122 281896
rect 399230 281808 399410 281896
rect 399518 281808 399698 281896
rect 399806 281808 399986 281896
rect 412286 281808 412466 281896
rect 412574 281808 412754 281896
rect 412862 281808 413042 281896
rect 413150 281808 413330 281896
rect 413438 281808 413618 281896
rect 413726 281808 413906 281896
rect 414014 281808 414194 281896
rect 414302 281808 414482 281896
rect 426782 281808 426962 281896
rect 427070 281808 427250 281896
rect 427358 281808 427538 281896
rect 427646 281808 427826 281896
rect 427934 281808 428114 281896
rect 428222 281808 428402 281896
rect 428510 281808 428690 281896
rect 428798 281808 428978 281896
rect 441278 281808 441458 281896
rect 441566 281808 441746 281896
rect 441854 281808 442034 281896
rect 442142 281808 442322 281896
rect 442430 281808 442610 281896
rect 442718 281808 442898 281896
rect 443006 281808 443186 281896
rect 443294 281808 443474 281896
rect 455774 281808 455954 281896
rect 456062 281808 456242 281896
rect 456350 281808 456530 281896
rect 456638 281808 456818 281896
rect 456926 281808 457106 281896
rect 457214 281808 457394 281896
rect 457502 281808 457682 281896
rect 457790 281808 457970 281896
rect 180350 281592 180530 281680
rect 180638 281592 180818 281680
rect 180926 281592 181106 281680
rect 181214 281592 181394 281680
rect 181502 281592 181682 281680
rect 181790 281592 181970 281680
rect 182078 281592 182258 281680
rect 182366 281592 182546 281680
rect 194846 281592 195026 281680
rect 195134 281592 195314 281680
rect 195422 281592 195602 281680
rect 195710 281592 195890 281680
rect 195998 281592 196178 281680
rect 196286 281592 196466 281680
rect 196574 281592 196754 281680
rect 196862 281592 197042 281680
rect 209342 281592 209522 281680
rect 209630 281592 209810 281680
rect 209918 281592 210098 281680
rect 210206 281592 210386 281680
rect 210494 281592 210674 281680
rect 210782 281592 210962 281680
rect 211070 281592 211250 281680
rect 211358 281592 211538 281680
rect 223838 281592 224018 281680
rect 224126 281592 224306 281680
rect 224414 281592 224594 281680
rect 224702 281592 224882 281680
rect 224990 281592 225170 281680
rect 225278 281592 225458 281680
rect 225566 281592 225746 281680
rect 225854 281592 226034 281680
rect 238334 281592 238514 281680
rect 238622 281592 238802 281680
rect 238910 281592 239090 281680
rect 239198 281592 239378 281680
rect 239486 281592 239666 281680
rect 239774 281592 239954 281680
rect 240062 281592 240242 281680
rect 240350 281592 240530 281680
rect 252830 281592 253010 281680
rect 253118 281592 253298 281680
rect 253406 281592 253586 281680
rect 253694 281592 253874 281680
rect 253982 281592 254162 281680
rect 254270 281592 254450 281680
rect 254558 281592 254738 281680
rect 254846 281592 255026 281680
rect 267326 281592 267506 281680
rect 267614 281592 267794 281680
rect 267902 281592 268082 281680
rect 268190 281592 268370 281680
rect 268478 281592 268658 281680
rect 268766 281592 268946 281680
rect 269054 281592 269234 281680
rect 269342 281592 269522 281680
rect 281822 281592 282002 281680
rect 282110 281592 282290 281680
rect 282398 281592 282578 281680
rect 282686 281592 282866 281680
rect 282974 281592 283154 281680
rect 283262 281592 283442 281680
rect 283550 281592 283730 281680
rect 283838 281592 284018 281680
rect 296318 281592 296498 281680
rect 296606 281592 296786 281680
rect 296894 281592 297074 281680
rect 297182 281592 297362 281680
rect 297470 281592 297650 281680
rect 297758 281592 297938 281680
rect 298046 281592 298226 281680
rect 298334 281592 298514 281680
rect 310814 281592 310994 281680
rect 311102 281592 311282 281680
rect 311390 281592 311570 281680
rect 311678 281592 311858 281680
rect 311966 281592 312146 281680
rect 312254 281592 312434 281680
rect 312542 281592 312722 281680
rect 312830 281592 313010 281680
rect 325310 281592 325490 281680
rect 325598 281592 325778 281680
rect 325886 281592 326066 281680
rect 326174 281592 326354 281680
rect 326462 281592 326642 281680
rect 326750 281592 326930 281680
rect 327038 281592 327218 281680
rect 327326 281592 327506 281680
rect 339806 281592 339986 281680
rect 340094 281592 340274 281680
rect 340382 281592 340562 281680
rect 340670 281592 340850 281680
rect 340958 281592 341138 281680
rect 341246 281592 341426 281680
rect 341534 281592 341714 281680
rect 341822 281592 342002 281680
rect 354302 281592 354482 281680
rect 354590 281592 354770 281680
rect 354878 281592 355058 281680
rect 355166 281592 355346 281680
rect 355454 281592 355634 281680
rect 355742 281592 355922 281680
rect 356030 281592 356210 281680
rect 356318 281592 356498 281680
rect 368798 281592 368978 281680
rect 369086 281592 369266 281680
rect 369374 281592 369554 281680
rect 369662 281592 369842 281680
rect 369950 281592 370130 281680
rect 370238 281592 370418 281680
rect 370526 281592 370706 281680
rect 370814 281592 370994 281680
rect 383294 281592 383474 281680
rect 383582 281592 383762 281680
rect 383870 281592 384050 281680
rect 384158 281592 384338 281680
rect 384446 281592 384626 281680
rect 384734 281592 384914 281680
rect 385022 281592 385202 281680
rect 385310 281592 385490 281680
rect 397790 281592 397970 281680
rect 398078 281592 398258 281680
rect 398366 281592 398546 281680
rect 398654 281592 398834 281680
rect 398942 281592 399122 281680
rect 399230 281592 399410 281680
rect 399518 281592 399698 281680
rect 399806 281592 399986 281680
rect 412286 281592 412466 281680
rect 412574 281592 412754 281680
rect 412862 281592 413042 281680
rect 413150 281592 413330 281680
rect 413438 281592 413618 281680
rect 413726 281592 413906 281680
rect 414014 281592 414194 281680
rect 414302 281592 414482 281680
rect 426782 281592 426962 281680
rect 427070 281592 427250 281680
rect 427358 281592 427538 281680
rect 427646 281592 427826 281680
rect 427934 281592 428114 281680
rect 428222 281592 428402 281680
rect 428510 281592 428690 281680
rect 428798 281592 428978 281680
rect 441278 281592 441458 281680
rect 441566 281592 441746 281680
rect 441854 281592 442034 281680
rect 442142 281592 442322 281680
rect 442430 281592 442610 281680
rect 442718 281592 442898 281680
rect 443006 281592 443186 281680
rect 443294 281592 443474 281680
rect 455774 281592 455954 281680
rect 456062 281592 456242 281680
rect 456350 281592 456530 281680
rect 456638 281592 456818 281680
rect 456926 281592 457106 281680
rect 457214 281592 457394 281680
rect 457502 281592 457682 281680
rect 457790 281592 457970 281680
rect 180350 281116 180530 281204
rect 180638 281116 180818 281204
rect 180926 281116 181106 281204
rect 181214 281116 181394 281204
rect 181502 281116 181682 281204
rect 181790 281116 181970 281204
rect 182078 281116 182258 281204
rect 182366 281116 182546 281204
rect 194846 281116 195026 281204
rect 195134 281116 195314 281204
rect 195422 281116 195602 281204
rect 195710 281116 195890 281204
rect 195998 281116 196178 281204
rect 196286 281116 196466 281204
rect 196574 281116 196754 281204
rect 196862 281116 197042 281204
rect 209342 281116 209522 281204
rect 209630 281116 209810 281204
rect 209918 281116 210098 281204
rect 210206 281116 210386 281204
rect 210494 281116 210674 281204
rect 210782 281116 210962 281204
rect 211070 281116 211250 281204
rect 211358 281116 211538 281204
rect 223838 281116 224018 281204
rect 224126 281116 224306 281204
rect 224414 281116 224594 281204
rect 224702 281116 224882 281204
rect 224990 281116 225170 281204
rect 225278 281116 225458 281204
rect 225566 281116 225746 281204
rect 225854 281116 226034 281204
rect 238334 281116 238514 281204
rect 238622 281116 238802 281204
rect 238910 281116 239090 281204
rect 239198 281116 239378 281204
rect 239486 281116 239666 281204
rect 239774 281116 239954 281204
rect 240062 281116 240242 281204
rect 240350 281116 240530 281204
rect 252830 281116 253010 281204
rect 253118 281116 253298 281204
rect 253406 281116 253586 281204
rect 253694 281116 253874 281204
rect 253982 281116 254162 281204
rect 254270 281116 254450 281204
rect 254558 281116 254738 281204
rect 254846 281116 255026 281204
rect 267326 281116 267506 281204
rect 267614 281116 267794 281204
rect 267902 281116 268082 281204
rect 268190 281116 268370 281204
rect 268478 281116 268658 281204
rect 268766 281116 268946 281204
rect 269054 281116 269234 281204
rect 269342 281116 269522 281204
rect 281822 281116 282002 281204
rect 282110 281116 282290 281204
rect 282398 281116 282578 281204
rect 282686 281116 282866 281204
rect 282974 281116 283154 281204
rect 283262 281116 283442 281204
rect 283550 281116 283730 281204
rect 283838 281116 284018 281204
rect 296318 281116 296498 281204
rect 296606 281116 296786 281204
rect 296894 281116 297074 281204
rect 297182 281116 297362 281204
rect 297470 281116 297650 281204
rect 297758 281116 297938 281204
rect 298046 281116 298226 281204
rect 298334 281116 298514 281204
rect 310814 281116 310994 281204
rect 311102 281116 311282 281204
rect 311390 281116 311570 281204
rect 311678 281116 311858 281204
rect 311966 281116 312146 281204
rect 312254 281116 312434 281204
rect 312542 281116 312722 281204
rect 312830 281116 313010 281204
rect 325310 281116 325490 281204
rect 325598 281116 325778 281204
rect 325886 281116 326066 281204
rect 326174 281116 326354 281204
rect 326462 281116 326642 281204
rect 326750 281116 326930 281204
rect 327038 281116 327218 281204
rect 327326 281116 327506 281204
rect 339806 281116 339986 281204
rect 340094 281116 340274 281204
rect 340382 281116 340562 281204
rect 340670 281116 340850 281204
rect 340958 281116 341138 281204
rect 341246 281116 341426 281204
rect 341534 281116 341714 281204
rect 341822 281116 342002 281204
rect 354302 281116 354482 281204
rect 354590 281116 354770 281204
rect 354878 281116 355058 281204
rect 355166 281116 355346 281204
rect 355454 281116 355634 281204
rect 355742 281116 355922 281204
rect 356030 281116 356210 281204
rect 356318 281116 356498 281204
rect 368798 281116 368978 281204
rect 369086 281116 369266 281204
rect 369374 281116 369554 281204
rect 369662 281116 369842 281204
rect 369950 281116 370130 281204
rect 370238 281116 370418 281204
rect 370526 281116 370706 281204
rect 370814 281116 370994 281204
rect 383294 281116 383474 281204
rect 383582 281116 383762 281204
rect 383870 281116 384050 281204
rect 384158 281116 384338 281204
rect 384446 281116 384626 281204
rect 384734 281116 384914 281204
rect 385022 281116 385202 281204
rect 385310 281116 385490 281204
rect 397790 281116 397970 281204
rect 398078 281116 398258 281204
rect 398366 281116 398546 281204
rect 398654 281116 398834 281204
rect 398942 281116 399122 281204
rect 399230 281116 399410 281204
rect 399518 281116 399698 281204
rect 399806 281116 399986 281204
rect 412286 281116 412466 281204
rect 412574 281116 412754 281204
rect 412862 281116 413042 281204
rect 413150 281116 413330 281204
rect 413438 281116 413618 281204
rect 413726 281116 413906 281204
rect 414014 281116 414194 281204
rect 414302 281116 414482 281204
rect 426782 281116 426962 281204
rect 427070 281116 427250 281204
rect 427358 281116 427538 281204
rect 427646 281116 427826 281204
rect 427934 281116 428114 281204
rect 428222 281116 428402 281204
rect 428510 281116 428690 281204
rect 428798 281116 428978 281204
rect 441278 281116 441458 281204
rect 441566 281116 441746 281204
rect 441854 281116 442034 281204
rect 442142 281116 442322 281204
rect 442430 281116 442610 281204
rect 442718 281116 442898 281204
rect 443006 281116 443186 281204
rect 443294 281116 443474 281204
rect 455774 281116 455954 281204
rect 456062 281116 456242 281204
rect 456350 281116 456530 281204
rect 456638 281116 456818 281204
rect 456926 281116 457106 281204
rect 457214 281116 457394 281204
rect 457502 281116 457682 281204
rect 457790 281116 457970 281204
rect 180350 280900 180530 280988
rect 180638 280900 180818 280988
rect 180926 280900 181106 280988
rect 181214 280900 181394 280988
rect 181502 280900 181682 280988
rect 181790 280900 181970 280988
rect 182078 280900 182258 280988
rect 182366 280900 182546 280988
rect 194846 280900 195026 280988
rect 195134 280900 195314 280988
rect 195422 280900 195602 280988
rect 195710 280900 195890 280988
rect 195998 280900 196178 280988
rect 196286 280900 196466 280988
rect 196574 280900 196754 280988
rect 196862 280900 197042 280988
rect 209342 280900 209522 280988
rect 209630 280900 209810 280988
rect 209918 280900 210098 280988
rect 210206 280900 210386 280988
rect 210494 280900 210674 280988
rect 210782 280900 210962 280988
rect 211070 280900 211250 280988
rect 211358 280900 211538 280988
rect 223838 280900 224018 280988
rect 224126 280900 224306 280988
rect 224414 280900 224594 280988
rect 224702 280900 224882 280988
rect 224990 280900 225170 280988
rect 225278 280900 225458 280988
rect 225566 280900 225746 280988
rect 225854 280900 226034 280988
rect 238334 280900 238514 280988
rect 238622 280900 238802 280988
rect 238910 280900 239090 280988
rect 239198 280900 239378 280988
rect 239486 280900 239666 280988
rect 239774 280900 239954 280988
rect 240062 280900 240242 280988
rect 240350 280900 240530 280988
rect 252830 280900 253010 280988
rect 253118 280900 253298 280988
rect 253406 280900 253586 280988
rect 253694 280900 253874 280988
rect 253982 280900 254162 280988
rect 254270 280900 254450 280988
rect 254558 280900 254738 280988
rect 254846 280900 255026 280988
rect 267326 280900 267506 280988
rect 267614 280900 267794 280988
rect 267902 280900 268082 280988
rect 268190 280900 268370 280988
rect 268478 280900 268658 280988
rect 268766 280900 268946 280988
rect 269054 280900 269234 280988
rect 269342 280900 269522 280988
rect 281822 280900 282002 280988
rect 282110 280900 282290 280988
rect 282398 280900 282578 280988
rect 282686 280900 282866 280988
rect 282974 280900 283154 280988
rect 283262 280900 283442 280988
rect 283550 280900 283730 280988
rect 283838 280900 284018 280988
rect 296318 280900 296498 280988
rect 296606 280900 296786 280988
rect 296894 280900 297074 280988
rect 297182 280900 297362 280988
rect 297470 280900 297650 280988
rect 297758 280900 297938 280988
rect 298046 280900 298226 280988
rect 298334 280900 298514 280988
rect 310814 280900 310994 280988
rect 311102 280900 311282 280988
rect 311390 280900 311570 280988
rect 311678 280900 311858 280988
rect 311966 280900 312146 280988
rect 312254 280900 312434 280988
rect 312542 280900 312722 280988
rect 312830 280900 313010 280988
rect 325310 280900 325490 280988
rect 325598 280900 325778 280988
rect 325886 280900 326066 280988
rect 326174 280900 326354 280988
rect 326462 280900 326642 280988
rect 326750 280900 326930 280988
rect 327038 280900 327218 280988
rect 327326 280900 327506 280988
rect 339806 280900 339986 280988
rect 340094 280900 340274 280988
rect 340382 280900 340562 280988
rect 340670 280900 340850 280988
rect 340958 280900 341138 280988
rect 341246 280900 341426 280988
rect 341534 280900 341714 280988
rect 341822 280900 342002 280988
rect 354302 280900 354482 280988
rect 354590 280900 354770 280988
rect 354878 280900 355058 280988
rect 355166 280900 355346 280988
rect 355454 280900 355634 280988
rect 355742 280900 355922 280988
rect 356030 280900 356210 280988
rect 356318 280900 356498 280988
rect 368798 280900 368978 280988
rect 369086 280900 369266 280988
rect 369374 280900 369554 280988
rect 369662 280900 369842 280988
rect 369950 280900 370130 280988
rect 370238 280900 370418 280988
rect 370526 280900 370706 280988
rect 370814 280900 370994 280988
rect 383294 280900 383474 280988
rect 383582 280900 383762 280988
rect 383870 280900 384050 280988
rect 384158 280900 384338 280988
rect 384446 280900 384626 280988
rect 384734 280900 384914 280988
rect 385022 280900 385202 280988
rect 385310 280900 385490 280988
rect 397790 280900 397970 280988
rect 398078 280900 398258 280988
rect 398366 280900 398546 280988
rect 398654 280900 398834 280988
rect 398942 280900 399122 280988
rect 399230 280900 399410 280988
rect 399518 280900 399698 280988
rect 399806 280900 399986 280988
rect 412286 280900 412466 280988
rect 412574 280900 412754 280988
rect 412862 280900 413042 280988
rect 413150 280900 413330 280988
rect 413438 280900 413618 280988
rect 413726 280900 413906 280988
rect 414014 280900 414194 280988
rect 414302 280900 414482 280988
rect 426782 280900 426962 280988
rect 427070 280900 427250 280988
rect 427358 280900 427538 280988
rect 427646 280900 427826 280988
rect 427934 280900 428114 280988
rect 428222 280900 428402 280988
rect 428510 280900 428690 280988
rect 428798 280900 428978 280988
rect 441278 280900 441458 280988
rect 441566 280900 441746 280988
rect 441854 280900 442034 280988
rect 442142 280900 442322 280988
rect 442430 280900 442610 280988
rect 442718 280900 442898 280988
rect 443006 280900 443186 280988
rect 443294 280900 443474 280988
rect 455774 280900 455954 280988
rect 456062 280900 456242 280988
rect 456350 280900 456530 280988
rect 456638 280900 456818 280988
rect 456926 280900 457106 280988
rect 457214 280900 457394 280988
rect 457502 280900 457682 280988
rect 457790 280900 457970 280988
rect 180350 266748 180530 266836
rect 180638 266748 180818 266836
rect 180926 266748 181106 266836
rect 181214 266748 181394 266836
rect 181502 266748 181682 266836
rect 181790 266748 181970 266836
rect 182078 266748 182258 266836
rect 182366 266748 182546 266836
rect 194846 266748 195026 266836
rect 195134 266748 195314 266836
rect 195422 266748 195602 266836
rect 195710 266748 195890 266836
rect 195998 266748 196178 266836
rect 196286 266748 196466 266836
rect 196574 266748 196754 266836
rect 196862 266748 197042 266836
rect 209342 266748 209522 266836
rect 209630 266748 209810 266836
rect 209918 266748 210098 266836
rect 210206 266748 210386 266836
rect 210494 266748 210674 266836
rect 210782 266748 210962 266836
rect 211070 266748 211250 266836
rect 211358 266748 211538 266836
rect 223838 266748 224018 266836
rect 224126 266748 224306 266836
rect 224414 266748 224594 266836
rect 224702 266748 224882 266836
rect 224990 266748 225170 266836
rect 225278 266748 225458 266836
rect 225566 266748 225746 266836
rect 225854 266748 226034 266836
rect 238334 266748 238514 266836
rect 238622 266748 238802 266836
rect 238910 266748 239090 266836
rect 239198 266748 239378 266836
rect 239486 266748 239666 266836
rect 239774 266748 239954 266836
rect 240062 266748 240242 266836
rect 240350 266748 240530 266836
rect 252830 266748 253010 266836
rect 253118 266748 253298 266836
rect 253406 266748 253586 266836
rect 253694 266748 253874 266836
rect 253982 266748 254162 266836
rect 254270 266748 254450 266836
rect 254558 266748 254738 266836
rect 254846 266748 255026 266836
rect 267326 266748 267506 266836
rect 267614 266748 267794 266836
rect 267902 266748 268082 266836
rect 268190 266748 268370 266836
rect 268478 266748 268658 266836
rect 268766 266748 268946 266836
rect 269054 266748 269234 266836
rect 269342 266748 269522 266836
rect 281822 266748 282002 266836
rect 282110 266748 282290 266836
rect 282398 266748 282578 266836
rect 282686 266748 282866 266836
rect 282974 266748 283154 266836
rect 283262 266748 283442 266836
rect 283550 266748 283730 266836
rect 283838 266748 284018 266836
rect 296318 266748 296498 266836
rect 296606 266748 296786 266836
rect 296894 266748 297074 266836
rect 297182 266748 297362 266836
rect 297470 266748 297650 266836
rect 297758 266748 297938 266836
rect 298046 266748 298226 266836
rect 298334 266748 298514 266836
rect 310814 266748 310994 266836
rect 311102 266748 311282 266836
rect 311390 266748 311570 266836
rect 311678 266748 311858 266836
rect 311966 266748 312146 266836
rect 312254 266748 312434 266836
rect 312542 266748 312722 266836
rect 312830 266748 313010 266836
rect 325310 266748 325490 266836
rect 325598 266748 325778 266836
rect 325886 266748 326066 266836
rect 326174 266748 326354 266836
rect 326462 266748 326642 266836
rect 326750 266748 326930 266836
rect 327038 266748 327218 266836
rect 327326 266748 327506 266836
rect 339806 266748 339986 266836
rect 340094 266748 340274 266836
rect 340382 266748 340562 266836
rect 340670 266748 340850 266836
rect 340958 266748 341138 266836
rect 341246 266748 341426 266836
rect 341534 266748 341714 266836
rect 341822 266748 342002 266836
rect 354302 266748 354482 266836
rect 354590 266748 354770 266836
rect 354878 266748 355058 266836
rect 355166 266748 355346 266836
rect 355454 266748 355634 266836
rect 355742 266748 355922 266836
rect 356030 266748 356210 266836
rect 356318 266748 356498 266836
rect 368798 266748 368978 266836
rect 369086 266748 369266 266836
rect 369374 266748 369554 266836
rect 369662 266748 369842 266836
rect 369950 266748 370130 266836
rect 370238 266748 370418 266836
rect 370526 266748 370706 266836
rect 370814 266748 370994 266836
rect 383294 266748 383474 266836
rect 383582 266748 383762 266836
rect 383870 266748 384050 266836
rect 384158 266748 384338 266836
rect 384446 266748 384626 266836
rect 384734 266748 384914 266836
rect 385022 266748 385202 266836
rect 385310 266748 385490 266836
rect 397790 266748 397970 266836
rect 398078 266748 398258 266836
rect 398366 266748 398546 266836
rect 398654 266748 398834 266836
rect 398942 266748 399122 266836
rect 399230 266748 399410 266836
rect 399518 266748 399698 266836
rect 399806 266748 399986 266836
rect 412286 266748 412466 266836
rect 412574 266748 412754 266836
rect 412862 266748 413042 266836
rect 413150 266748 413330 266836
rect 413438 266748 413618 266836
rect 413726 266748 413906 266836
rect 414014 266748 414194 266836
rect 414302 266748 414482 266836
rect 426782 266748 426962 266836
rect 427070 266748 427250 266836
rect 427358 266748 427538 266836
rect 427646 266748 427826 266836
rect 427934 266748 428114 266836
rect 428222 266748 428402 266836
rect 428510 266748 428690 266836
rect 428798 266748 428978 266836
rect 441278 266748 441458 266836
rect 441566 266748 441746 266836
rect 441854 266748 442034 266836
rect 442142 266748 442322 266836
rect 442430 266748 442610 266836
rect 442718 266748 442898 266836
rect 443006 266748 443186 266836
rect 443294 266748 443474 266836
rect 455774 266748 455954 266836
rect 456062 266748 456242 266836
rect 456350 266748 456530 266836
rect 456638 266748 456818 266836
rect 456926 266748 457106 266836
rect 457214 266748 457394 266836
rect 457502 266748 457682 266836
rect 457790 266748 457970 266836
rect 180350 266532 180530 266620
rect 180638 266532 180818 266620
rect 180926 266532 181106 266620
rect 181214 266532 181394 266620
rect 181502 266532 181682 266620
rect 181790 266532 181970 266620
rect 182078 266532 182258 266620
rect 182366 266532 182546 266620
rect 194846 266532 195026 266620
rect 195134 266532 195314 266620
rect 195422 266532 195602 266620
rect 195710 266532 195890 266620
rect 195998 266532 196178 266620
rect 196286 266532 196466 266620
rect 196574 266532 196754 266620
rect 196862 266532 197042 266620
rect 209342 266532 209522 266620
rect 209630 266532 209810 266620
rect 209918 266532 210098 266620
rect 210206 266532 210386 266620
rect 210494 266532 210674 266620
rect 210782 266532 210962 266620
rect 211070 266532 211250 266620
rect 211358 266532 211538 266620
rect 223838 266532 224018 266620
rect 224126 266532 224306 266620
rect 224414 266532 224594 266620
rect 224702 266532 224882 266620
rect 224990 266532 225170 266620
rect 225278 266532 225458 266620
rect 225566 266532 225746 266620
rect 225854 266532 226034 266620
rect 238334 266532 238514 266620
rect 238622 266532 238802 266620
rect 238910 266532 239090 266620
rect 239198 266532 239378 266620
rect 239486 266532 239666 266620
rect 239774 266532 239954 266620
rect 240062 266532 240242 266620
rect 240350 266532 240530 266620
rect 252830 266532 253010 266620
rect 253118 266532 253298 266620
rect 253406 266532 253586 266620
rect 253694 266532 253874 266620
rect 253982 266532 254162 266620
rect 254270 266532 254450 266620
rect 254558 266532 254738 266620
rect 254846 266532 255026 266620
rect 267326 266532 267506 266620
rect 267614 266532 267794 266620
rect 267902 266532 268082 266620
rect 268190 266532 268370 266620
rect 268478 266532 268658 266620
rect 268766 266532 268946 266620
rect 269054 266532 269234 266620
rect 269342 266532 269522 266620
rect 281822 266532 282002 266620
rect 282110 266532 282290 266620
rect 282398 266532 282578 266620
rect 282686 266532 282866 266620
rect 282974 266532 283154 266620
rect 283262 266532 283442 266620
rect 283550 266532 283730 266620
rect 283838 266532 284018 266620
rect 296318 266532 296498 266620
rect 296606 266532 296786 266620
rect 296894 266532 297074 266620
rect 297182 266532 297362 266620
rect 297470 266532 297650 266620
rect 297758 266532 297938 266620
rect 298046 266532 298226 266620
rect 298334 266532 298514 266620
rect 310814 266532 310994 266620
rect 311102 266532 311282 266620
rect 311390 266532 311570 266620
rect 311678 266532 311858 266620
rect 311966 266532 312146 266620
rect 312254 266532 312434 266620
rect 312542 266532 312722 266620
rect 312830 266532 313010 266620
rect 325310 266532 325490 266620
rect 325598 266532 325778 266620
rect 325886 266532 326066 266620
rect 326174 266532 326354 266620
rect 326462 266532 326642 266620
rect 326750 266532 326930 266620
rect 327038 266532 327218 266620
rect 327326 266532 327506 266620
rect 339806 266532 339986 266620
rect 340094 266532 340274 266620
rect 340382 266532 340562 266620
rect 340670 266532 340850 266620
rect 340958 266532 341138 266620
rect 341246 266532 341426 266620
rect 341534 266532 341714 266620
rect 341822 266532 342002 266620
rect 354302 266532 354482 266620
rect 354590 266532 354770 266620
rect 354878 266532 355058 266620
rect 355166 266532 355346 266620
rect 355454 266532 355634 266620
rect 355742 266532 355922 266620
rect 356030 266532 356210 266620
rect 356318 266532 356498 266620
rect 368798 266532 368978 266620
rect 369086 266532 369266 266620
rect 369374 266532 369554 266620
rect 369662 266532 369842 266620
rect 369950 266532 370130 266620
rect 370238 266532 370418 266620
rect 370526 266532 370706 266620
rect 370814 266532 370994 266620
rect 383294 266532 383474 266620
rect 383582 266532 383762 266620
rect 383870 266532 384050 266620
rect 384158 266532 384338 266620
rect 384446 266532 384626 266620
rect 384734 266532 384914 266620
rect 385022 266532 385202 266620
rect 385310 266532 385490 266620
rect 397790 266532 397970 266620
rect 398078 266532 398258 266620
rect 398366 266532 398546 266620
rect 398654 266532 398834 266620
rect 398942 266532 399122 266620
rect 399230 266532 399410 266620
rect 399518 266532 399698 266620
rect 399806 266532 399986 266620
rect 412286 266532 412466 266620
rect 412574 266532 412754 266620
rect 412862 266532 413042 266620
rect 413150 266532 413330 266620
rect 413438 266532 413618 266620
rect 413726 266532 413906 266620
rect 414014 266532 414194 266620
rect 414302 266532 414482 266620
rect 426782 266532 426962 266620
rect 427070 266532 427250 266620
rect 427358 266532 427538 266620
rect 427646 266532 427826 266620
rect 427934 266532 428114 266620
rect 428222 266532 428402 266620
rect 428510 266532 428690 266620
rect 428798 266532 428978 266620
rect 441278 266532 441458 266620
rect 441566 266532 441746 266620
rect 441854 266532 442034 266620
rect 442142 266532 442322 266620
rect 442430 266532 442610 266620
rect 442718 266532 442898 266620
rect 443006 266532 443186 266620
rect 443294 266532 443474 266620
rect 455774 266532 455954 266620
rect 456062 266532 456242 266620
rect 456350 266532 456530 266620
rect 456638 266532 456818 266620
rect 456926 266532 457106 266620
rect 457214 266532 457394 266620
rect 457502 266532 457682 266620
rect 457790 266532 457970 266620
rect 180350 266056 180530 266144
rect 180638 266056 180818 266144
rect 180926 266056 181106 266144
rect 181214 266056 181394 266144
rect 181502 266056 181682 266144
rect 181790 266056 181970 266144
rect 182078 266056 182258 266144
rect 182366 266056 182546 266144
rect 194846 266056 195026 266144
rect 195134 266056 195314 266144
rect 195422 266056 195602 266144
rect 195710 266056 195890 266144
rect 195998 266056 196178 266144
rect 196286 266056 196466 266144
rect 196574 266056 196754 266144
rect 196862 266056 197042 266144
rect 209342 266056 209522 266144
rect 209630 266056 209810 266144
rect 209918 266056 210098 266144
rect 210206 266056 210386 266144
rect 210494 266056 210674 266144
rect 210782 266056 210962 266144
rect 211070 266056 211250 266144
rect 211358 266056 211538 266144
rect 223838 266056 224018 266144
rect 224126 266056 224306 266144
rect 224414 266056 224594 266144
rect 224702 266056 224882 266144
rect 224990 266056 225170 266144
rect 225278 266056 225458 266144
rect 225566 266056 225746 266144
rect 225854 266056 226034 266144
rect 238334 266056 238514 266144
rect 238622 266056 238802 266144
rect 238910 266056 239090 266144
rect 239198 266056 239378 266144
rect 239486 266056 239666 266144
rect 239774 266056 239954 266144
rect 240062 266056 240242 266144
rect 240350 266056 240530 266144
rect 252830 266056 253010 266144
rect 253118 266056 253298 266144
rect 253406 266056 253586 266144
rect 253694 266056 253874 266144
rect 253982 266056 254162 266144
rect 254270 266056 254450 266144
rect 254558 266056 254738 266144
rect 254846 266056 255026 266144
rect 267326 266056 267506 266144
rect 267614 266056 267794 266144
rect 267902 266056 268082 266144
rect 268190 266056 268370 266144
rect 268478 266056 268658 266144
rect 268766 266056 268946 266144
rect 269054 266056 269234 266144
rect 269342 266056 269522 266144
rect 281822 266056 282002 266144
rect 282110 266056 282290 266144
rect 282398 266056 282578 266144
rect 282686 266056 282866 266144
rect 282974 266056 283154 266144
rect 283262 266056 283442 266144
rect 283550 266056 283730 266144
rect 283838 266056 284018 266144
rect 296318 266056 296498 266144
rect 296606 266056 296786 266144
rect 296894 266056 297074 266144
rect 297182 266056 297362 266144
rect 297470 266056 297650 266144
rect 297758 266056 297938 266144
rect 298046 266056 298226 266144
rect 298334 266056 298514 266144
rect 310814 266056 310994 266144
rect 311102 266056 311282 266144
rect 311390 266056 311570 266144
rect 311678 266056 311858 266144
rect 311966 266056 312146 266144
rect 312254 266056 312434 266144
rect 312542 266056 312722 266144
rect 312830 266056 313010 266144
rect 325310 266056 325490 266144
rect 325598 266056 325778 266144
rect 325886 266056 326066 266144
rect 326174 266056 326354 266144
rect 326462 266056 326642 266144
rect 326750 266056 326930 266144
rect 327038 266056 327218 266144
rect 327326 266056 327506 266144
rect 339806 266056 339986 266144
rect 340094 266056 340274 266144
rect 340382 266056 340562 266144
rect 340670 266056 340850 266144
rect 340958 266056 341138 266144
rect 341246 266056 341426 266144
rect 341534 266056 341714 266144
rect 341822 266056 342002 266144
rect 354302 266056 354482 266144
rect 354590 266056 354770 266144
rect 354878 266056 355058 266144
rect 355166 266056 355346 266144
rect 355454 266056 355634 266144
rect 355742 266056 355922 266144
rect 356030 266056 356210 266144
rect 356318 266056 356498 266144
rect 368798 266056 368978 266144
rect 369086 266056 369266 266144
rect 369374 266056 369554 266144
rect 369662 266056 369842 266144
rect 369950 266056 370130 266144
rect 370238 266056 370418 266144
rect 370526 266056 370706 266144
rect 370814 266056 370994 266144
rect 383294 266056 383474 266144
rect 383582 266056 383762 266144
rect 383870 266056 384050 266144
rect 384158 266056 384338 266144
rect 384446 266056 384626 266144
rect 384734 266056 384914 266144
rect 385022 266056 385202 266144
rect 385310 266056 385490 266144
rect 397790 266056 397970 266144
rect 398078 266056 398258 266144
rect 398366 266056 398546 266144
rect 398654 266056 398834 266144
rect 398942 266056 399122 266144
rect 399230 266056 399410 266144
rect 399518 266056 399698 266144
rect 399806 266056 399986 266144
rect 412286 266056 412466 266144
rect 412574 266056 412754 266144
rect 412862 266056 413042 266144
rect 413150 266056 413330 266144
rect 413438 266056 413618 266144
rect 413726 266056 413906 266144
rect 414014 266056 414194 266144
rect 414302 266056 414482 266144
rect 426782 266056 426962 266144
rect 427070 266056 427250 266144
rect 427358 266056 427538 266144
rect 427646 266056 427826 266144
rect 427934 266056 428114 266144
rect 428222 266056 428402 266144
rect 428510 266056 428690 266144
rect 428798 266056 428978 266144
rect 441278 266056 441458 266144
rect 441566 266056 441746 266144
rect 441854 266056 442034 266144
rect 442142 266056 442322 266144
rect 442430 266056 442610 266144
rect 442718 266056 442898 266144
rect 443006 266056 443186 266144
rect 443294 266056 443474 266144
rect 455774 266056 455954 266144
rect 456062 266056 456242 266144
rect 456350 266056 456530 266144
rect 456638 266056 456818 266144
rect 456926 266056 457106 266144
rect 457214 266056 457394 266144
rect 457502 266056 457682 266144
rect 457790 266056 457970 266144
rect 180350 265840 180530 265928
rect 180638 265840 180818 265928
rect 180926 265840 181106 265928
rect 181214 265840 181394 265928
rect 181502 265840 181682 265928
rect 181790 265840 181970 265928
rect 182078 265840 182258 265928
rect 182366 265840 182546 265928
rect 194846 265840 195026 265928
rect 195134 265840 195314 265928
rect 195422 265840 195602 265928
rect 195710 265840 195890 265928
rect 195998 265840 196178 265928
rect 196286 265840 196466 265928
rect 196574 265840 196754 265928
rect 196862 265840 197042 265928
rect 209342 265840 209522 265928
rect 209630 265840 209810 265928
rect 209918 265840 210098 265928
rect 210206 265840 210386 265928
rect 210494 265840 210674 265928
rect 210782 265840 210962 265928
rect 211070 265840 211250 265928
rect 211358 265840 211538 265928
rect 223838 265840 224018 265928
rect 224126 265840 224306 265928
rect 224414 265840 224594 265928
rect 224702 265840 224882 265928
rect 224990 265840 225170 265928
rect 225278 265840 225458 265928
rect 225566 265840 225746 265928
rect 225854 265840 226034 265928
rect 238334 265840 238514 265928
rect 238622 265840 238802 265928
rect 238910 265840 239090 265928
rect 239198 265840 239378 265928
rect 239486 265840 239666 265928
rect 239774 265840 239954 265928
rect 240062 265840 240242 265928
rect 240350 265840 240530 265928
rect 252830 265840 253010 265928
rect 253118 265840 253298 265928
rect 253406 265840 253586 265928
rect 253694 265840 253874 265928
rect 253982 265840 254162 265928
rect 254270 265840 254450 265928
rect 254558 265840 254738 265928
rect 254846 265840 255026 265928
rect 267326 265840 267506 265928
rect 267614 265840 267794 265928
rect 267902 265840 268082 265928
rect 268190 265840 268370 265928
rect 268478 265840 268658 265928
rect 268766 265840 268946 265928
rect 269054 265840 269234 265928
rect 269342 265840 269522 265928
rect 281822 265840 282002 265928
rect 282110 265840 282290 265928
rect 282398 265840 282578 265928
rect 282686 265840 282866 265928
rect 282974 265840 283154 265928
rect 283262 265840 283442 265928
rect 283550 265840 283730 265928
rect 283838 265840 284018 265928
rect 296318 265840 296498 265928
rect 296606 265840 296786 265928
rect 296894 265840 297074 265928
rect 297182 265840 297362 265928
rect 297470 265840 297650 265928
rect 297758 265840 297938 265928
rect 298046 265840 298226 265928
rect 298334 265840 298514 265928
rect 310814 265840 310994 265928
rect 311102 265840 311282 265928
rect 311390 265840 311570 265928
rect 311678 265840 311858 265928
rect 311966 265840 312146 265928
rect 312254 265840 312434 265928
rect 312542 265840 312722 265928
rect 312830 265840 313010 265928
rect 325310 265840 325490 265928
rect 325598 265840 325778 265928
rect 325886 265840 326066 265928
rect 326174 265840 326354 265928
rect 326462 265840 326642 265928
rect 326750 265840 326930 265928
rect 327038 265840 327218 265928
rect 327326 265840 327506 265928
rect 339806 265840 339986 265928
rect 340094 265840 340274 265928
rect 340382 265840 340562 265928
rect 340670 265840 340850 265928
rect 340958 265840 341138 265928
rect 341246 265840 341426 265928
rect 341534 265840 341714 265928
rect 341822 265840 342002 265928
rect 354302 265840 354482 265928
rect 354590 265840 354770 265928
rect 354878 265840 355058 265928
rect 355166 265840 355346 265928
rect 355454 265840 355634 265928
rect 355742 265840 355922 265928
rect 356030 265840 356210 265928
rect 356318 265840 356498 265928
rect 368798 265840 368978 265928
rect 369086 265840 369266 265928
rect 369374 265840 369554 265928
rect 369662 265840 369842 265928
rect 369950 265840 370130 265928
rect 370238 265840 370418 265928
rect 370526 265840 370706 265928
rect 370814 265840 370994 265928
rect 383294 265840 383474 265928
rect 383582 265840 383762 265928
rect 383870 265840 384050 265928
rect 384158 265840 384338 265928
rect 384446 265840 384626 265928
rect 384734 265840 384914 265928
rect 385022 265840 385202 265928
rect 385310 265840 385490 265928
rect 397790 265840 397970 265928
rect 398078 265840 398258 265928
rect 398366 265840 398546 265928
rect 398654 265840 398834 265928
rect 398942 265840 399122 265928
rect 399230 265840 399410 265928
rect 399518 265840 399698 265928
rect 399806 265840 399986 265928
rect 412286 265840 412466 265928
rect 412574 265840 412754 265928
rect 412862 265840 413042 265928
rect 413150 265840 413330 265928
rect 413438 265840 413618 265928
rect 413726 265840 413906 265928
rect 414014 265840 414194 265928
rect 414302 265840 414482 265928
rect 426782 265840 426962 265928
rect 427070 265840 427250 265928
rect 427358 265840 427538 265928
rect 427646 265840 427826 265928
rect 427934 265840 428114 265928
rect 428222 265840 428402 265928
rect 428510 265840 428690 265928
rect 428798 265840 428978 265928
rect 441278 265840 441458 265928
rect 441566 265840 441746 265928
rect 441854 265840 442034 265928
rect 442142 265840 442322 265928
rect 442430 265840 442610 265928
rect 442718 265840 442898 265928
rect 443006 265840 443186 265928
rect 443294 265840 443474 265928
rect 455774 265840 455954 265928
rect 456062 265840 456242 265928
rect 456350 265840 456530 265928
rect 456638 265840 456818 265928
rect 456926 265840 457106 265928
rect 457214 265840 457394 265928
rect 457502 265840 457682 265928
rect 457790 265840 457970 265928
rect 180350 251688 180530 251776
rect 180638 251688 180818 251776
rect 180926 251688 181106 251776
rect 181214 251688 181394 251776
rect 181502 251688 181682 251776
rect 181790 251688 181970 251776
rect 182078 251688 182258 251776
rect 182366 251688 182546 251776
rect 194846 251688 195026 251776
rect 195134 251688 195314 251776
rect 195422 251688 195602 251776
rect 195710 251688 195890 251776
rect 195998 251688 196178 251776
rect 196286 251688 196466 251776
rect 196574 251688 196754 251776
rect 196862 251688 197042 251776
rect 209342 251688 209522 251776
rect 209630 251688 209810 251776
rect 209918 251688 210098 251776
rect 210206 251688 210386 251776
rect 210494 251688 210674 251776
rect 210782 251688 210962 251776
rect 211070 251688 211250 251776
rect 211358 251688 211538 251776
rect 223838 251688 224018 251776
rect 224126 251688 224306 251776
rect 224414 251688 224594 251776
rect 224702 251688 224882 251776
rect 224990 251688 225170 251776
rect 225278 251688 225458 251776
rect 225566 251688 225746 251776
rect 225854 251688 226034 251776
rect 238334 251688 238514 251776
rect 238622 251688 238802 251776
rect 238910 251688 239090 251776
rect 239198 251688 239378 251776
rect 239486 251688 239666 251776
rect 239774 251688 239954 251776
rect 240062 251688 240242 251776
rect 240350 251688 240530 251776
rect 252830 251688 253010 251776
rect 253118 251688 253298 251776
rect 253406 251688 253586 251776
rect 253694 251688 253874 251776
rect 253982 251688 254162 251776
rect 254270 251688 254450 251776
rect 254558 251688 254738 251776
rect 254846 251688 255026 251776
rect 267326 251688 267506 251776
rect 267614 251688 267794 251776
rect 267902 251688 268082 251776
rect 268190 251688 268370 251776
rect 268478 251688 268658 251776
rect 268766 251688 268946 251776
rect 269054 251688 269234 251776
rect 269342 251688 269522 251776
rect 281822 251688 282002 251776
rect 282110 251688 282290 251776
rect 282398 251688 282578 251776
rect 282686 251688 282866 251776
rect 282974 251688 283154 251776
rect 283262 251688 283442 251776
rect 283550 251688 283730 251776
rect 283838 251688 284018 251776
rect 296318 251688 296498 251776
rect 296606 251688 296786 251776
rect 296894 251688 297074 251776
rect 297182 251688 297362 251776
rect 297470 251688 297650 251776
rect 297758 251688 297938 251776
rect 298046 251688 298226 251776
rect 298334 251688 298514 251776
rect 310814 251688 310994 251776
rect 311102 251688 311282 251776
rect 311390 251688 311570 251776
rect 311678 251688 311858 251776
rect 311966 251688 312146 251776
rect 312254 251688 312434 251776
rect 312542 251688 312722 251776
rect 312830 251688 313010 251776
rect 325310 251688 325490 251776
rect 325598 251688 325778 251776
rect 325886 251688 326066 251776
rect 326174 251688 326354 251776
rect 326462 251688 326642 251776
rect 326750 251688 326930 251776
rect 327038 251688 327218 251776
rect 327326 251688 327506 251776
rect 339806 251688 339986 251776
rect 340094 251688 340274 251776
rect 340382 251688 340562 251776
rect 340670 251688 340850 251776
rect 340958 251688 341138 251776
rect 341246 251688 341426 251776
rect 341534 251688 341714 251776
rect 341822 251688 342002 251776
rect 354302 251688 354482 251776
rect 354590 251688 354770 251776
rect 354878 251688 355058 251776
rect 355166 251688 355346 251776
rect 355454 251688 355634 251776
rect 355742 251688 355922 251776
rect 356030 251688 356210 251776
rect 356318 251688 356498 251776
rect 368798 251688 368978 251776
rect 369086 251688 369266 251776
rect 369374 251688 369554 251776
rect 369662 251688 369842 251776
rect 369950 251688 370130 251776
rect 370238 251688 370418 251776
rect 370526 251688 370706 251776
rect 370814 251688 370994 251776
rect 383294 251688 383474 251776
rect 383582 251688 383762 251776
rect 383870 251688 384050 251776
rect 384158 251688 384338 251776
rect 384446 251688 384626 251776
rect 384734 251688 384914 251776
rect 385022 251688 385202 251776
rect 385310 251688 385490 251776
rect 397790 251688 397970 251776
rect 398078 251688 398258 251776
rect 398366 251688 398546 251776
rect 398654 251688 398834 251776
rect 398942 251688 399122 251776
rect 399230 251688 399410 251776
rect 399518 251688 399698 251776
rect 399806 251688 399986 251776
rect 412286 251688 412466 251776
rect 412574 251688 412754 251776
rect 412862 251688 413042 251776
rect 413150 251688 413330 251776
rect 413438 251688 413618 251776
rect 413726 251688 413906 251776
rect 414014 251688 414194 251776
rect 414302 251688 414482 251776
rect 426782 251688 426962 251776
rect 427070 251688 427250 251776
rect 427358 251688 427538 251776
rect 427646 251688 427826 251776
rect 427934 251688 428114 251776
rect 428222 251688 428402 251776
rect 428510 251688 428690 251776
rect 428798 251688 428978 251776
rect 441278 251688 441458 251776
rect 441566 251688 441746 251776
rect 441854 251688 442034 251776
rect 442142 251688 442322 251776
rect 442430 251688 442610 251776
rect 442718 251688 442898 251776
rect 443006 251688 443186 251776
rect 443294 251688 443474 251776
rect 455774 251688 455954 251776
rect 456062 251688 456242 251776
rect 456350 251688 456530 251776
rect 456638 251688 456818 251776
rect 456926 251688 457106 251776
rect 457214 251688 457394 251776
rect 457502 251688 457682 251776
rect 457790 251688 457970 251776
rect 180350 251472 180530 251560
rect 180638 251472 180818 251560
rect 180926 251472 181106 251560
rect 181214 251472 181394 251560
rect 181502 251472 181682 251560
rect 181790 251472 181970 251560
rect 182078 251472 182258 251560
rect 182366 251472 182546 251560
rect 194846 251472 195026 251560
rect 195134 251472 195314 251560
rect 195422 251472 195602 251560
rect 195710 251472 195890 251560
rect 195998 251472 196178 251560
rect 196286 251472 196466 251560
rect 196574 251472 196754 251560
rect 196862 251472 197042 251560
rect 209342 251472 209522 251560
rect 209630 251472 209810 251560
rect 209918 251472 210098 251560
rect 210206 251472 210386 251560
rect 210494 251472 210674 251560
rect 210782 251472 210962 251560
rect 211070 251472 211250 251560
rect 211358 251472 211538 251560
rect 223838 251472 224018 251560
rect 224126 251472 224306 251560
rect 224414 251472 224594 251560
rect 224702 251472 224882 251560
rect 224990 251472 225170 251560
rect 225278 251472 225458 251560
rect 225566 251472 225746 251560
rect 225854 251472 226034 251560
rect 238334 251472 238514 251560
rect 238622 251472 238802 251560
rect 238910 251472 239090 251560
rect 239198 251472 239378 251560
rect 239486 251472 239666 251560
rect 239774 251472 239954 251560
rect 240062 251472 240242 251560
rect 240350 251472 240530 251560
rect 252830 251472 253010 251560
rect 253118 251472 253298 251560
rect 253406 251472 253586 251560
rect 253694 251472 253874 251560
rect 253982 251472 254162 251560
rect 254270 251472 254450 251560
rect 254558 251472 254738 251560
rect 254846 251472 255026 251560
rect 267326 251472 267506 251560
rect 267614 251472 267794 251560
rect 267902 251472 268082 251560
rect 268190 251472 268370 251560
rect 268478 251472 268658 251560
rect 268766 251472 268946 251560
rect 269054 251472 269234 251560
rect 269342 251472 269522 251560
rect 281822 251472 282002 251560
rect 282110 251472 282290 251560
rect 282398 251472 282578 251560
rect 282686 251472 282866 251560
rect 282974 251472 283154 251560
rect 283262 251472 283442 251560
rect 283550 251472 283730 251560
rect 283838 251472 284018 251560
rect 296318 251472 296498 251560
rect 296606 251472 296786 251560
rect 296894 251472 297074 251560
rect 297182 251472 297362 251560
rect 297470 251472 297650 251560
rect 297758 251472 297938 251560
rect 298046 251472 298226 251560
rect 298334 251472 298514 251560
rect 310814 251472 310994 251560
rect 311102 251472 311282 251560
rect 311390 251472 311570 251560
rect 311678 251472 311858 251560
rect 311966 251472 312146 251560
rect 312254 251472 312434 251560
rect 312542 251472 312722 251560
rect 312830 251472 313010 251560
rect 325310 251472 325490 251560
rect 325598 251472 325778 251560
rect 325886 251472 326066 251560
rect 326174 251472 326354 251560
rect 326462 251472 326642 251560
rect 326750 251472 326930 251560
rect 327038 251472 327218 251560
rect 327326 251472 327506 251560
rect 339806 251472 339986 251560
rect 340094 251472 340274 251560
rect 340382 251472 340562 251560
rect 340670 251472 340850 251560
rect 340958 251472 341138 251560
rect 341246 251472 341426 251560
rect 341534 251472 341714 251560
rect 341822 251472 342002 251560
rect 354302 251472 354482 251560
rect 354590 251472 354770 251560
rect 354878 251472 355058 251560
rect 355166 251472 355346 251560
rect 355454 251472 355634 251560
rect 355742 251472 355922 251560
rect 356030 251472 356210 251560
rect 356318 251472 356498 251560
rect 368798 251472 368978 251560
rect 369086 251472 369266 251560
rect 369374 251472 369554 251560
rect 369662 251472 369842 251560
rect 369950 251472 370130 251560
rect 370238 251472 370418 251560
rect 370526 251472 370706 251560
rect 370814 251472 370994 251560
rect 383294 251472 383474 251560
rect 383582 251472 383762 251560
rect 383870 251472 384050 251560
rect 384158 251472 384338 251560
rect 384446 251472 384626 251560
rect 384734 251472 384914 251560
rect 385022 251472 385202 251560
rect 385310 251472 385490 251560
rect 397790 251472 397970 251560
rect 398078 251472 398258 251560
rect 398366 251472 398546 251560
rect 398654 251472 398834 251560
rect 398942 251472 399122 251560
rect 399230 251472 399410 251560
rect 399518 251472 399698 251560
rect 399806 251472 399986 251560
rect 412286 251472 412466 251560
rect 412574 251472 412754 251560
rect 412862 251472 413042 251560
rect 413150 251472 413330 251560
rect 413438 251472 413618 251560
rect 413726 251472 413906 251560
rect 414014 251472 414194 251560
rect 414302 251472 414482 251560
rect 426782 251472 426962 251560
rect 427070 251472 427250 251560
rect 427358 251472 427538 251560
rect 427646 251472 427826 251560
rect 427934 251472 428114 251560
rect 428222 251472 428402 251560
rect 428510 251472 428690 251560
rect 428798 251472 428978 251560
rect 441278 251472 441458 251560
rect 441566 251472 441746 251560
rect 441854 251472 442034 251560
rect 442142 251472 442322 251560
rect 442430 251472 442610 251560
rect 442718 251472 442898 251560
rect 443006 251472 443186 251560
rect 443294 251472 443474 251560
rect 455774 251472 455954 251560
rect 456062 251472 456242 251560
rect 456350 251472 456530 251560
rect 456638 251472 456818 251560
rect 456926 251472 457106 251560
rect 457214 251472 457394 251560
rect 457502 251472 457682 251560
rect 457790 251472 457970 251560
rect 180350 250996 180530 251084
rect 180638 250996 180818 251084
rect 180926 250996 181106 251084
rect 181214 250996 181394 251084
rect 181502 250996 181682 251084
rect 181790 250996 181970 251084
rect 182078 250996 182258 251084
rect 182366 250996 182546 251084
rect 194846 250996 195026 251084
rect 195134 250996 195314 251084
rect 195422 250996 195602 251084
rect 195710 250996 195890 251084
rect 195998 250996 196178 251084
rect 196286 250996 196466 251084
rect 196574 250996 196754 251084
rect 196862 250996 197042 251084
rect 209342 250996 209522 251084
rect 209630 250996 209810 251084
rect 209918 250996 210098 251084
rect 210206 250996 210386 251084
rect 210494 250996 210674 251084
rect 210782 250996 210962 251084
rect 211070 250996 211250 251084
rect 211358 250996 211538 251084
rect 223838 250996 224018 251084
rect 224126 250996 224306 251084
rect 224414 250996 224594 251084
rect 224702 250996 224882 251084
rect 224990 250996 225170 251084
rect 225278 250996 225458 251084
rect 225566 250996 225746 251084
rect 225854 250996 226034 251084
rect 238334 250996 238514 251084
rect 238622 250996 238802 251084
rect 238910 250996 239090 251084
rect 239198 250996 239378 251084
rect 239486 250996 239666 251084
rect 239774 250996 239954 251084
rect 240062 250996 240242 251084
rect 240350 250996 240530 251084
rect 252830 250996 253010 251084
rect 253118 250996 253298 251084
rect 253406 250996 253586 251084
rect 253694 250996 253874 251084
rect 253982 250996 254162 251084
rect 254270 250996 254450 251084
rect 254558 250996 254738 251084
rect 254846 250996 255026 251084
rect 267326 250996 267506 251084
rect 267614 250996 267794 251084
rect 267902 250996 268082 251084
rect 268190 250996 268370 251084
rect 268478 250996 268658 251084
rect 268766 250996 268946 251084
rect 269054 250996 269234 251084
rect 269342 250996 269522 251084
rect 281822 250996 282002 251084
rect 282110 250996 282290 251084
rect 282398 250996 282578 251084
rect 282686 250996 282866 251084
rect 282974 250996 283154 251084
rect 283262 250996 283442 251084
rect 283550 250996 283730 251084
rect 283838 250996 284018 251084
rect 296318 250996 296498 251084
rect 296606 250996 296786 251084
rect 296894 250996 297074 251084
rect 297182 250996 297362 251084
rect 297470 250996 297650 251084
rect 297758 250996 297938 251084
rect 298046 250996 298226 251084
rect 298334 250996 298514 251084
rect 310814 250996 310994 251084
rect 311102 250996 311282 251084
rect 311390 250996 311570 251084
rect 311678 250996 311858 251084
rect 311966 250996 312146 251084
rect 312254 250996 312434 251084
rect 312542 250996 312722 251084
rect 312830 250996 313010 251084
rect 325310 250996 325490 251084
rect 325598 250996 325778 251084
rect 325886 250996 326066 251084
rect 326174 250996 326354 251084
rect 326462 250996 326642 251084
rect 326750 250996 326930 251084
rect 327038 250996 327218 251084
rect 327326 250996 327506 251084
rect 339806 250996 339986 251084
rect 340094 250996 340274 251084
rect 340382 250996 340562 251084
rect 340670 250996 340850 251084
rect 340958 250996 341138 251084
rect 341246 250996 341426 251084
rect 341534 250996 341714 251084
rect 341822 250996 342002 251084
rect 354302 250996 354482 251084
rect 354590 250996 354770 251084
rect 354878 250996 355058 251084
rect 355166 250996 355346 251084
rect 355454 250996 355634 251084
rect 355742 250996 355922 251084
rect 356030 250996 356210 251084
rect 356318 250996 356498 251084
rect 368798 250996 368978 251084
rect 369086 250996 369266 251084
rect 369374 250996 369554 251084
rect 369662 250996 369842 251084
rect 369950 250996 370130 251084
rect 370238 250996 370418 251084
rect 370526 250996 370706 251084
rect 370814 250996 370994 251084
rect 383294 250996 383474 251084
rect 383582 250996 383762 251084
rect 383870 250996 384050 251084
rect 384158 250996 384338 251084
rect 384446 250996 384626 251084
rect 384734 250996 384914 251084
rect 385022 250996 385202 251084
rect 385310 250996 385490 251084
rect 397790 250996 397970 251084
rect 398078 250996 398258 251084
rect 398366 250996 398546 251084
rect 398654 250996 398834 251084
rect 398942 250996 399122 251084
rect 399230 250996 399410 251084
rect 399518 250996 399698 251084
rect 399806 250996 399986 251084
rect 412286 250996 412466 251084
rect 412574 250996 412754 251084
rect 412862 250996 413042 251084
rect 413150 250996 413330 251084
rect 413438 250996 413618 251084
rect 413726 250996 413906 251084
rect 414014 250996 414194 251084
rect 414302 250996 414482 251084
rect 426782 250996 426962 251084
rect 427070 250996 427250 251084
rect 427358 250996 427538 251084
rect 427646 250996 427826 251084
rect 427934 250996 428114 251084
rect 428222 250996 428402 251084
rect 428510 250996 428690 251084
rect 428798 250996 428978 251084
rect 441278 250996 441458 251084
rect 441566 250996 441746 251084
rect 441854 250996 442034 251084
rect 442142 250996 442322 251084
rect 442430 250996 442610 251084
rect 442718 250996 442898 251084
rect 443006 250996 443186 251084
rect 443294 250996 443474 251084
rect 455774 250996 455954 251084
rect 456062 250996 456242 251084
rect 456350 250996 456530 251084
rect 456638 250996 456818 251084
rect 456926 250996 457106 251084
rect 457214 250996 457394 251084
rect 457502 250996 457682 251084
rect 457790 250996 457970 251084
rect 180350 250780 180530 250868
rect 180638 250780 180818 250868
rect 180926 250780 181106 250868
rect 181214 250780 181394 250868
rect 181502 250780 181682 250868
rect 181790 250780 181970 250868
rect 182078 250780 182258 250868
rect 182366 250780 182546 250868
rect 194846 250780 195026 250868
rect 195134 250780 195314 250868
rect 195422 250780 195602 250868
rect 195710 250780 195890 250868
rect 195998 250780 196178 250868
rect 196286 250780 196466 250868
rect 196574 250780 196754 250868
rect 196862 250780 197042 250868
rect 209342 250780 209522 250868
rect 209630 250780 209810 250868
rect 209918 250780 210098 250868
rect 210206 250780 210386 250868
rect 210494 250780 210674 250868
rect 210782 250780 210962 250868
rect 211070 250780 211250 250868
rect 211358 250780 211538 250868
rect 223838 250780 224018 250868
rect 224126 250780 224306 250868
rect 224414 250780 224594 250868
rect 224702 250780 224882 250868
rect 224990 250780 225170 250868
rect 225278 250780 225458 250868
rect 225566 250780 225746 250868
rect 225854 250780 226034 250868
rect 238334 250780 238514 250868
rect 238622 250780 238802 250868
rect 238910 250780 239090 250868
rect 239198 250780 239378 250868
rect 239486 250780 239666 250868
rect 239774 250780 239954 250868
rect 240062 250780 240242 250868
rect 240350 250780 240530 250868
rect 252830 250780 253010 250868
rect 253118 250780 253298 250868
rect 253406 250780 253586 250868
rect 253694 250780 253874 250868
rect 253982 250780 254162 250868
rect 254270 250780 254450 250868
rect 254558 250780 254738 250868
rect 254846 250780 255026 250868
rect 267326 250780 267506 250868
rect 267614 250780 267794 250868
rect 267902 250780 268082 250868
rect 268190 250780 268370 250868
rect 268478 250780 268658 250868
rect 268766 250780 268946 250868
rect 269054 250780 269234 250868
rect 269342 250780 269522 250868
rect 281822 250780 282002 250868
rect 282110 250780 282290 250868
rect 282398 250780 282578 250868
rect 282686 250780 282866 250868
rect 282974 250780 283154 250868
rect 283262 250780 283442 250868
rect 283550 250780 283730 250868
rect 283838 250780 284018 250868
rect 296318 250780 296498 250868
rect 296606 250780 296786 250868
rect 296894 250780 297074 250868
rect 297182 250780 297362 250868
rect 297470 250780 297650 250868
rect 297758 250780 297938 250868
rect 298046 250780 298226 250868
rect 298334 250780 298514 250868
rect 310814 250780 310994 250868
rect 311102 250780 311282 250868
rect 311390 250780 311570 250868
rect 311678 250780 311858 250868
rect 311966 250780 312146 250868
rect 312254 250780 312434 250868
rect 312542 250780 312722 250868
rect 312830 250780 313010 250868
rect 325310 250780 325490 250868
rect 325598 250780 325778 250868
rect 325886 250780 326066 250868
rect 326174 250780 326354 250868
rect 326462 250780 326642 250868
rect 326750 250780 326930 250868
rect 327038 250780 327218 250868
rect 327326 250780 327506 250868
rect 339806 250780 339986 250868
rect 340094 250780 340274 250868
rect 340382 250780 340562 250868
rect 340670 250780 340850 250868
rect 340958 250780 341138 250868
rect 341246 250780 341426 250868
rect 341534 250780 341714 250868
rect 341822 250780 342002 250868
rect 354302 250780 354482 250868
rect 354590 250780 354770 250868
rect 354878 250780 355058 250868
rect 355166 250780 355346 250868
rect 355454 250780 355634 250868
rect 355742 250780 355922 250868
rect 356030 250780 356210 250868
rect 356318 250780 356498 250868
rect 368798 250780 368978 250868
rect 369086 250780 369266 250868
rect 369374 250780 369554 250868
rect 369662 250780 369842 250868
rect 369950 250780 370130 250868
rect 370238 250780 370418 250868
rect 370526 250780 370706 250868
rect 370814 250780 370994 250868
rect 383294 250780 383474 250868
rect 383582 250780 383762 250868
rect 383870 250780 384050 250868
rect 384158 250780 384338 250868
rect 384446 250780 384626 250868
rect 384734 250780 384914 250868
rect 385022 250780 385202 250868
rect 385310 250780 385490 250868
rect 397790 250780 397970 250868
rect 398078 250780 398258 250868
rect 398366 250780 398546 250868
rect 398654 250780 398834 250868
rect 398942 250780 399122 250868
rect 399230 250780 399410 250868
rect 399518 250780 399698 250868
rect 399806 250780 399986 250868
rect 412286 250780 412466 250868
rect 412574 250780 412754 250868
rect 412862 250780 413042 250868
rect 413150 250780 413330 250868
rect 413438 250780 413618 250868
rect 413726 250780 413906 250868
rect 414014 250780 414194 250868
rect 414302 250780 414482 250868
rect 426782 250780 426962 250868
rect 427070 250780 427250 250868
rect 427358 250780 427538 250868
rect 427646 250780 427826 250868
rect 427934 250780 428114 250868
rect 428222 250780 428402 250868
rect 428510 250780 428690 250868
rect 428798 250780 428978 250868
rect 441278 250780 441458 250868
rect 441566 250780 441746 250868
rect 441854 250780 442034 250868
rect 442142 250780 442322 250868
rect 442430 250780 442610 250868
rect 442718 250780 442898 250868
rect 443006 250780 443186 250868
rect 443294 250780 443474 250868
rect 455774 250780 455954 250868
rect 456062 250780 456242 250868
rect 456350 250780 456530 250868
rect 456638 250780 456818 250868
rect 456926 250780 457106 250868
rect 457214 250780 457394 250868
rect 457502 250780 457682 250868
rect 457790 250780 457970 250868
rect 180350 236628 180530 236716
rect 180638 236628 180818 236716
rect 180926 236628 181106 236716
rect 181214 236628 181394 236716
rect 181502 236628 181682 236716
rect 181790 236628 181970 236716
rect 182078 236628 182258 236716
rect 182366 236628 182546 236716
rect 194846 236628 195026 236716
rect 195134 236628 195314 236716
rect 195422 236628 195602 236716
rect 195710 236628 195890 236716
rect 195998 236628 196178 236716
rect 196286 236628 196466 236716
rect 196574 236628 196754 236716
rect 196862 236628 197042 236716
rect 209342 236628 209522 236716
rect 209630 236628 209810 236716
rect 209918 236628 210098 236716
rect 210206 236628 210386 236716
rect 210494 236628 210674 236716
rect 210782 236628 210962 236716
rect 211070 236628 211250 236716
rect 211358 236628 211538 236716
rect 223838 236628 224018 236716
rect 224126 236628 224306 236716
rect 224414 236628 224594 236716
rect 224702 236628 224882 236716
rect 224990 236628 225170 236716
rect 225278 236628 225458 236716
rect 225566 236628 225746 236716
rect 225854 236628 226034 236716
rect 238334 236628 238514 236716
rect 238622 236628 238802 236716
rect 238910 236628 239090 236716
rect 239198 236628 239378 236716
rect 239486 236628 239666 236716
rect 239774 236628 239954 236716
rect 240062 236628 240242 236716
rect 240350 236628 240530 236716
rect 252830 236628 253010 236716
rect 253118 236628 253298 236716
rect 253406 236628 253586 236716
rect 253694 236628 253874 236716
rect 253982 236628 254162 236716
rect 254270 236628 254450 236716
rect 254558 236628 254738 236716
rect 254846 236628 255026 236716
rect 267326 236628 267506 236716
rect 267614 236628 267794 236716
rect 267902 236628 268082 236716
rect 268190 236628 268370 236716
rect 268478 236628 268658 236716
rect 268766 236628 268946 236716
rect 269054 236628 269234 236716
rect 269342 236628 269522 236716
rect 281822 236628 282002 236716
rect 282110 236628 282290 236716
rect 282398 236628 282578 236716
rect 282686 236628 282866 236716
rect 282974 236628 283154 236716
rect 283262 236628 283442 236716
rect 283550 236628 283730 236716
rect 283838 236628 284018 236716
rect 296318 236628 296498 236716
rect 296606 236628 296786 236716
rect 296894 236628 297074 236716
rect 297182 236628 297362 236716
rect 297470 236628 297650 236716
rect 297758 236628 297938 236716
rect 298046 236628 298226 236716
rect 298334 236628 298514 236716
rect 310814 236628 310994 236716
rect 311102 236628 311282 236716
rect 311390 236628 311570 236716
rect 311678 236628 311858 236716
rect 311966 236628 312146 236716
rect 312254 236628 312434 236716
rect 312542 236628 312722 236716
rect 312830 236628 313010 236716
rect 325310 236628 325490 236716
rect 325598 236628 325778 236716
rect 325886 236628 326066 236716
rect 326174 236628 326354 236716
rect 326462 236628 326642 236716
rect 326750 236628 326930 236716
rect 327038 236628 327218 236716
rect 327326 236628 327506 236716
rect 339806 236628 339986 236716
rect 340094 236628 340274 236716
rect 340382 236628 340562 236716
rect 340670 236628 340850 236716
rect 340958 236628 341138 236716
rect 341246 236628 341426 236716
rect 341534 236628 341714 236716
rect 341822 236628 342002 236716
rect 354302 236628 354482 236716
rect 354590 236628 354770 236716
rect 354878 236628 355058 236716
rect 355166 236628 355346 236716
rect 355454 236628 355634 236716
rect 355742 236628 355922 236716
rect 356030 236628 356210 236716
rect 356318 236628 356498 236716
rect 368798 236628 368978 236716
rect 369086 236628 369266 236716
rect 369374 236628 369554 236716
rect 369662 236628 369842 236716
rect 369950 236628 370130 236716
rect 370238 236628 370418 236716
rect 370526 236628 370706 236716
rect 370814 236628 370994 236716
rect 383294 236628 383474 236716
rect 383582 236628 383762 236716
rect 383870 236628 384050 236716
rect 384158 236628 384338 236716
rect 384446 236628 384626 236716
rect 384734 236628 384914 236716
rect 385022 236628 385202 236716
rect 385310 236628 385490 236716
rect 397790 236628 397970 236716
rect 398078 236628 398258 236716
rect 398366 236628 398546 236716
rect 398654 236628 398834 236716
rect 398942 236628 399122 236716
rect 399230 236628 399410 236716
rect 399518 236628 399698 236716
rect 399806 236628 399986 236716
rect 412286 236628 412466 236716
rect 412574 236628 412754 236716
rect 412862 236628 413042 236716
rect 413150 236628 413330 236716
rect 413438 236628 413618 236716
rect 413726 236628 413906 236716
rect 414014 236628 414194 236716
rect 414302 236628 414482 236716
rect 426782 236628 426962 236716
rect 427070 236628 427250 236716
rect 427358 236628 427538 236716
rect 427646 236628 427826 236716
rect 427934 236628 428114 236716
rect 428222 236628 428402 236716
rect 428510 236628 428690 236716
rect 428798 236628 428978 236716
rect 441278 236628 441458 236716
rect 441566 236628 441746 236716
rect 441854 236628 442034 236716
rect 442142 236628 442322 236716
rect 442430 236628 442610 236716
rect 442718 236628 442898 236716
rect 443006 236628 443186 236716
rect 443294 236628 443474 236716
rect 455774 236628 455954 236716
rect 456062 236628 456242 236716
rect 456350 236628 456530 236716
rect 456638 236628 456818 236716
rect 456926 236628 457106 236716
rect 457214 236628 457394 236716
rect 457502 236628 457682 236716
rect 457790 236628 457970 236716
rect 180350 236412 180530 236500
rect 180638 236412 180818 236500
rect 180926 236412 181106 236500
rect 181214 236412 181394 236500
rect 181502 236412 181682 236500
rect 181790 236412 181970 236500
rect 182078 236412 182258 236500
rect 182366 236412 182546 236500
rect 194846 236412 195026 236500
rect 195134 236412 195314 236500
rect 195422 236412 195602 236500
rect 195710 236412 195890 236500
rect 195998 236412 196178 236500
rect 196286 236412 196466 236500
rect 196574 236412 196754 236500
rect 196862 236412 197042 236500
rect 209342 236412 209522 236500
rect 209630 236412 209810 236500
rect 209918 236412 210098 236500
rect 210206 236412 210386 236500
rect 210494 236412 210674 236500
rect 210782 236412 210962 236500
rect 211070 236412 211250 236500
rect 211358 236412 211538 236500
rect 223838 236412 224018 236500
rect 224126 236412 224306 236500
rect 224414 236412 224594 236500
rect 224702 236412 224882 236500
rect 224990 236412 225170 236500
rect 225278 236412 225458 236500
rect 225566 236412 225746 236500
rect 225854 236412 226034 236500
rect 238334 236412 238514 236500
rect 238622 236412 238802 236500
rect 238910 236412 239090 236500
rect 239198 236412 239378 236500
rect 239486 236412 239666 236500
rect 239774 236412 239954 236500
rect 240062 236412 240242 236500
rect 240350 236412 240530 236500
rect 252830 236412 253010 236500
rect 253118 236412 253298 236500
rect 253406 236412 253586 236500
rect 253694 236412 253874 236500
rect 253982 236412 254162 236500
rect 254270 236412 254450 236500
rect 254558 236412 254738 236500
rect 254846 236412 255026 236500
rect 267326 236412 267506 236500
rect 267614 236412 267794 236500
rect 267902 236412 268082 236500
rect 268190 236412 268370 236500
rect 268478 236412 268658 236500
rect 268766 236412 268946 236500
rect 269054 236412 269234 236500
rect 269342 236412 269522 236500
rect 281822 236412 282002 236500
rect 282110 236412 282290 236500
rect 282398 236412 282578 236500
rect 282686 236412 282866 236500
rect 282974 236412 283154 236500
rect 283262 236412 283442 236500
rect 283550 236412 283730 236500
rect 283838 236412 284018 236500
rect 296318 236412 296498 236500
rect 296606 236412 296786 236500
rect 296894 236412 297074 236500
rect 297182 236412 297362 236500
rect 297470 236412 297650 236500
rect 297758 236412 297938 236500
rect 298046 236412 298226 236500
rect 298334 236412 298514 236500
rect 310814 236412 310994 236500
rect 311102 236412 311282 236500
rect 311390 236412 311570 236500
rect 311678 236412 311858 236500
rect 311966 236412 312146 236500
rect 312254 236412 312434 236500
rect 312542 236412 312722 236500
rect 312830 236412 313010 236500
rect 325310 236412 325490 236500
rect 325598 236412 325778 236500
rect 325886 236412 326066 236500
rect 326174 236412 326354 236500
rect 326462 236412 326642 236500
rect 326750 236412 326930 236500
rect 327038 236412 327218 236500
rect 327326 236412 327506 236500
rect 339806 236412 339986 236500
rect 340094 236412 340274 236500
rect 340382 236412 340562 236500
rect 340670 236412 340850 236500
rect 340958 236412 341138 236500
rect 341246 236412 341426 236500
rect 341534 236412 341714 236500
rect 341822 236412 342002 236500
rect 354302 236412 354482 236500
rect 354590 236412 354770 236500
rect 354878 236412 355058 236500
rect 355166 236412 355346 236500
rect 355454 236412 355634 236500
rect 355742 236412 355922 236500
rect 356030 236412 356210 236500
rect 356318 236412 356498 236500
rect 368798 236412 368978 236500
rect 369086 236412 369266 236500
rect 369374 236412 369554 236500
rect 369662 236412 369842 236500
rect 369950 236412 370130 236500
rect 370238 236412 370418 236500
rect 370526 236412 370706 236500
rect 370814 236412 370994 236500
rect 383294 236412 383474 236500
rect 383582 236412 383762 236500
rect 383870 236412 384050 236500
rect 384158 236412 384338 236500
rect 384446 236412 384626 236500
rect 384734 236412 384914 236500
rect 385022 236412 385202 236500
rect 385310 236412 385490 236500
rect 397790 236412 397970 236500
rect 398078 236412 398258 236500
rect 398366 236412 398546 236500
rect 398654 236412 398834 236500
rect 398942 236412 399122 236500
rect 399230 236412 399410 236500
rect 399518 236412 399698 236500
rect 399806 236412 399986 236500
rect 412286 236412 412466 236500
rect 412574 236412 412754 236500
rect 412862 236412 413042 236500
rect 413150 236412 413330 236500
rect 413438 236412 413618 236500
rect 413726 236412 413906 236500
rect 414014 236412 414194 236500
rect 414302 236412 414482 236500
rect 426782 236412 426962 236500
rect 427070 236412 427250 236500
rect 427358 236412 427538 236500
rect 427646 236412 427826 236500
rect 427934 236412 428114 236500
rect 428222 236412 428402 236500
rect 428510 236412 428690 236500
rect 428798 236412 428978 236500
rect 441278 236412 441458 236500
rect 441566 236412 441746 236500
rect 441854 236412 442034 236500
rect 442142 236412 442322 236500
rect 442430 236412 442610 236500
rect 442718 236412 442898 236500
rect 443006 236412 443186 236500
rect 443294 236412 443474 236500
rect 455774 236412 455954 236500
rect 456062 236412 456242 236500
rect 456350 236412 456530 236500
rect 456638 236412 456818 236500
rect 456926 236412 457106 236500
rect 457214 236412 457394 236500
rect 457502 236412 457682 236500
rect 457790 236412 457970 236500
rect 180350 235936 180530 236024
rect 180638 235936 180818 236024
rect 180926 235936 181106 236024
rect 181214 235936 181394 236024
rect 181502 235936 181682 236024
rect 181790 235936 181970 236024
rect 182078 235936 182258 236024
rect 182366 235936 182546 236024
rect 194846 235936 195026 236024
rect 195134 235936 195314 236024
rect 195422 235936 195602 236024
rect 195710 235936 195890 236024
rect 195998 235936 196178 236024
rect 196286 235936 196466 236024
rect 196574 235936 196754 236024
rect 196862 235936 197042 236024
rect 209342 235936 209522 236024
rect 209630 235936 209810 236024
rect 209918 235936 210098 236024
rect 210206 235936 210386 236024
rect 210494 235936 210674 236024
rect 210782 235936 210962 236024
rect 211070 235936 211250 236024
rect 211358 235936 211538 236024
rect 223838 235936 224018 236024
rect 224126 235936 224306 236024
rect 224414 235936 224594 236024
rect 224702 235936 224882 236024
rect 224990 235936 225170 236024
rect 225278 235936 225458 236024
rect 225566 235936 225746 236024
rect 225854 235936 226034 236024
rect 238334 235936 238514 236024
rect 238622 235936 238802 236024
rect 238910 235936 239090 236024
rect 239198 235936 239378 236024
rect 239486 235936 239666 236024
rect 239774 235936 239954 236024
rect 240062 235936 240242 236024
rect 240350 235936 240530 236024
rect 252830 235936 253010 236024
rect 253118 235936 253298 236024
rect 253406 235936 253586 236024
rect 253694 235936 253874 236024
rect 253982 235936 254162 236024
rect 254270 235936 254450 236024
rect 254558 235936 254738 236024
rect 254846 235936 255026 236024
rect 267326 235936 267506 236024
rect 267614 235936 267794 236024
rect 267902 235936 268082 236024
rect 268190 235936 268370 236024
rect 268478 235936 268658 236024
rect 268766 235936 268946 236024
rect 269054 235936 269234 236024
rect 269342 235936 269522 236024
rect 281822 235936 282002 236024
rect 282110 235936 282290 236024
rect 282398 235936 282578 236024
rect 282686 235936 282866 236024
rect 282974 235936 283154 236024
rect 283262 235936 283442 236024
rect 283550 235936 283730 236024
rect 283838 235936 284018 236024
rect 296318 235936 296498 236024
rect 296606 235936 296786 236024
rect 296894 235936 297074 236024
rect 297182 235936 297362 236024
rect 297470 235936 297650 236024
rect 297758 235936 297938 236024
rect 298046 235936 298226 236024
rect 298334 235936 298514 236024
rect 310814 235936 310994 236024
rect 311102 235936 311282 236024
rect 311390 235936 311570 236024
rect 311678 235936 311858 236024
rect 311966 235936 312146 236024
rect 312254 235936 312434 236024
rect 312542 235936 312722 236024
rect 312830 235936 313010 236024
rect 325310 235936 325490 236024
rect 325598 235936 325778 236024
rect 325886 235936 326066 236024
rect 326174 235936 326354 236024
rect 326462 235936 326642 236024
rect 326750 235936 326930 236024
rect 327038 235936 327218 236024
rect 327326 235936 327506 236024
rect 339806 235936 339986 236024
rect 340094 235936 340274 236024
rect 340382 235936 340562 236024
rect 340670 235936 340850 236024
rect 340958 235936 341138 236024
rect 341246 235936 341426 236024
rect 341534 235936 341714 236024
rect 341822 235936 342002 236024
rect 354302 235936 354482 236024
rect 354590 235936 354770 236024
rect 354878 235936 355058 236024
rect 355166 235936 355346 236024
rect 355454 235936 355634 236024
rect 355742 235936 355922 236024
rect 356030 235936 356210 236024
rect 356318 235936 356498 236024
rect 368798 235936 368978 236024
rect 369086 235936 369266 236024
rect 369374 235936 369554 236024
rect 369662 235936 369842 236024
rect 369950 235936 370130 236024
rect 370238 235936 370418 236024
rect 370526 235936 370706 236024
rect 370814 235936 370994 236024
rect 383294 235936 383474 236024
rect 383582 235936 383762 236024
rect 383870 235936 384050 236024
rect 384158 235936 384338 236024
rect 384446 235936 384626 236024
rect 384734 235936 384914 236024
rect 385022 235936 385202 236024
rect 385310 235936 385490 236024
rect 397790 235936 397970 236024
rect 398078 235936 398258 236024
rect 398366 235936 398546 236024
rect 398654 235936 398834 236024
rect 398942 235936 399122 236024
rect 399230 235936 399410 236024
rect 399518 235936 399698 236024
rect 399806 235936 399986 236024
rect 412286 235936 412466 236024
rect 412574 235936 412754 236024
rect 412862 235936 413042 236024
rect 413150 235936 413330 236024
rect 413438 235936 413618 236024
rect 413726 235936 413906 236024
rect 414014 235936 414194 236024
rect 414302 235936 414482 236024
rect 426782 235936 426962 236024
rect 427070 235936 427250 236024
rect 427358 235936 427538 236024
rect 427646 235936 427826 236024
rect 427934 235936 428114 236024
rect 428222 235936 428402 236024
rect 428510 235936 428690 236024
rect 428798 235936 428978 236024
rect 441278 235936 441458 236024
rect 441566 235936 441746 236024
rect 441854 235936 442034 236024
rect 442142 235936 442322 236024
rect 442430 235936 442610 236024
rect 442718 235936 442898 236024
rect 443006 235936 443186 236024
rect 443294 235936 443474 236024
rect 455774 235936 455954 236024
rect 456062 235936 456242 236024
rect 456350 235936 456530 236024
rect 456638 235936 456818 236024
rect 456926 235936 457106 236024
rect 457214 235936 457394 236024
rect 457502 235936 457682 236024
rect 457790 235936 457970 236024
rect 180350 235720 180530 235808
rect 180638 235720 180818 235808
rect 180926 235720 181106 235808
rect 181214 235720 181394 235808
rect 181502 235720 181682 235808
rect 181790 235720 181970 235808
rect 182078 235720 182258 235808
rect 182366 235720 182546 235808
rect 194846 235720 195026 235808
rect 195134 235720 195314 235808
rect 195422 235720 195602 235808
rect 195710 235720 195890 235808
rect 195998 235720 196178 235808
rect 196286 235720 196466 235808
rect 196574 235720 196754 235808
rect 196862 235720 197042 235808
rect 209342 235720 209522 235808
rect 209630 235720 209810 235808
rect 209918 235720 210098 235808
rect 210206 235720 210386 235808
rect 210494 235720 210674 235808
rect 210782 235720 210962 235808
rect 211070 235720 211250 235808
rect 211358 235720 211538 235808
rect 223838 235720 224018 235808
rect 224126 235720 224306 235808
rect 224414 235720 224594 235808
rect 224702 235720 224882 235808
rect 224990 235720 225170 235808
rect 225278 235720 225458 235808
rect 225566 235720 225746 235808
rect 225854 235720 226034 235808
rect 238334 235720 238514 235808
rect 238622 235720 238802 235808
rect 238910 235720 239090 235808
rect 239198 235720 239378 235808
rect 239486 235720 239666 235808
rect 239774 235720 239954 235808
rect 240062 235720 240242 235808
rect 240350 235720 240530 235808
rect 252830 235720 253010 235808
rect 253118 235720 253298 235808
rect 253406 235720 253586 235808
rect 253694 235720 253874 235808
rect 253982 235720 254162 235808
rect 254270 235720 254450 235808
rect 254558 235720 254738 235808
rect 254846 235720 255026 235808
rect 267326 235720 267506 235808
rect 267614 235720 267794 235808
rect 267902 235720 268082 235808
rect 268190 235720 268370 235808
rect 268478 235720 268658 235808
rect 268766 235720 268946 235808
rect 269054 235720 269234 235808
rect 269342 235720 269522 235808
rect 281822 235720 282002 235808
rect 282110 235720 282290 235808
rect 282398 235720 282578 235808
rect 282686 235720 282866 235808
rect 282974 235720 283154 235808
rect 283262 235720 283442 235808
rect 283550 235720 283730 235808
rect 283838 235720 284018 235808
rect 296318 235720 296498 235808
rect 296606 235720 296786 235808
rect 296894 235720 297074 235808
rect 297182 235720 297362 235808
rect 297470 235720 297650 235808
rect 297758 235720 297938 235808
rect 298046 235720 298226 235808
rect 298334 235720 298514 235808
rect 310814 235720 310994 235808
rect 311102 235720 311282 235808
rect 311390 235720 311570 235808
rect 311678 235720 311858 235808
rect 311966 235720 312146 235808
rect 312254 235720 312434 235808
rect 312542 235720 312722 235808
rect 312830 235720 313010 235808
rect 325310 235720 325490 235808
rect 325598 235720 325778 235808
rect 325886 235720 326066 235808
rect 326174 235720 326354 235808
rect 326462 235720 326642 235808
rect 326750 235720 326930 235808
rect 327038 235720 327218 235808
rect 327326 235720 327506 235808
rect 339806 235720 339986 235808
rect 340094 235720 340274 235808
rect 340382 235720 340562 235808
rect 340670 235720 340850 235808
rect 340958 235720 341138 235808
rect 341246 235720 341426 235808
rect 341534 235720 341714 235808
rect 341822 235720 342002 235808
rect 354302 235720 354482 235808
rect 354590 235720 354770 235808
rect 354878 235720 355058 235808
rect 355166 235720 355346 235808
rect 355454 235720 355634 235808
rect 355742 235720 355922 235808
rect 356030 235720 356210 235808
rect 356318 235720 356498 235808
rect 368798 235720 368978 235808
rect 369086 235720 369266 235808
rect 369374 235720 369554 235808
rect 369662 235720 369842 235808
rect 369950 235720 370130 235808
rect 370238 235720 370418 235808
rect 370526 235720 370706 235808
rect 370814 235720 370994 235808
rect 383294 235720 383474 235808
rect 383582 235720 383762 235808
rect 383870 235720 384050 235808
rect 384158 235720 384338 235808
rect 384446 235720 384626 235808
rect 384734 235720 384914 235808
rect 385022 235720 385202 235808
rect 385310 235720 385490 235808
rect 397790 235720 397970 235808
rect 398078 235720 398258 235808
rect 398366 235720 398546 235808
rect 398654 235720 398834 235808
rect 398942 235720 399122 235808
rect 399230 235720 399410 235808
rect 399518 235720 399698 235808
rect 399806 235720 399986 235808
rect 412286 235720 412466 235808
rect 412574 235720 412754 235808
rect 412862 235720 413042 235808
rect 413150 235720 413330 235808
rect 413438 235720 413618 235808
rect 413726 235720 413906 235808
rect 414014 235720 414194 235808
rect 414302 235720 414482 235808
rect 426782 235720 426962 235808
rect 427070 235720 427250 235808
rect 427358 235720 427538 235808
rect 427646 235720 427826 235808
rect 427934 235720 428114 235808
rect 428222 235720 428402 235808
rect 428510 235720 428690 235808
rect 428798 235720 428978 235808
rect 441278 235720 441458 235808
rect 441566 235720 441746 235808
rect 441854 235720 442034 235808
rect 442142 235720 442322 235808
rect 442430 235720 442610 235808
rect 442718 235720 442898 235808
rect 443006 235720 443186 235808
rect 443294 235720 443474 235808
rect 455774 235720 455954 235808
rect 456062 235720 456242 235808
rect 456350 235720 456530 235808
rect 456638 235720 456818 235808
rect 456926 235720 457106 235808
rect 457214 235720 457394 235808
rect 457502 235720 457682 235808
rect 457790 235720 457970 235808
rect 180350 221568 180530 221656
rect 180638 221568 180818 221656
rect 180926 221568 181106 221656
rect 181214 221568 181394 221656
rect 181502 221568 181682 221656
rect 181790 221568 181970 221656
rect 182078 221568 182258 221656
rect 182366 221568 182546 221656
rect 194846 221568 195026 221656
rect 195134 221568 195314 221656
rect 195422 221568 195602 221656
rect 195710 221568 195890 221656
rect 195998 221568 196178 221656
rect 196286 221568 196466 221656
rect 196574 221568 196754 221656
rect 196862 221568 197042 221656
rect 209342 221568 209522 221656
rect 209630 221568 209810 221656
rect 209918 221568 210098 221656
rect 210206 221568 210386 221656
rect 210494 221568 210674 221656
rect 210782 221568 210962 221656
rect 211070 221568 211250 221656
rect 211358 221568 211538 221656
rect 223838 221568 224018 221656
rect 224126 221568 224306 221656
rect 224414 221568 224594 221656
rect 224702 221568 224882 221656
rect 224990 221568 225170 221656
rect 225278 221568 225458 221656
rect 225566 221568 225746 221656
rect 225854 221568 226034 221656
rect 238334 221568 238514 221656
rect 238622 221568 238802 221656
rect 238910 221568 239090 221656
rect 239198 221568 239378 221656
rect 239486 221568 239666 221656
rect 239774 221568 239954 221656
rect 240062 221568 240242 221656
rect 240350 221568 240530 221656
rect 252830 221568 253010 221656
rect 253118 221568 253298 221656
rect 253406 221568 253586 221656
rect 253694 221568 253874 221656
rect 253982 221568 254162 221656
rect 254270 221568 254450 221656
rect 254558 221568 254738 221656
rect 254846 221568 255026 221656
rect 267326 221568 267506 221656
rect 267614 221568 267794 221656
rect 267902 221568 268082 221656
rect 268190 221568 268370 221656
rect 268478 221568 268658 221656
rect 268766 221568 268946 221656
rect 269054 221568 269234 221656
rect 269342 221568 269522 221656
rect 281822 221568 282002 221656
rect 282110 221568 282290 221656
rect 282398 221568 282578 221656
rect 282686 221568 282866 221656
rect 282974 221568 283154 221656
rect 283262 221568 283442 221656
rect 283550 221568 283730 221656
rect 283838 221568 284018 221656
rect 296318 221568 296498 221656
rect 296606 221568 296786 221656
rect 296894 221568 297074 221656
rect 297182 221568 297362 221656
rect 297470 221568 297650 221656
rect 297758 221568 297938 221656
rect 298046 221568 298226 221656
rect 298334 221568 298514 221656
rect 310814 221568 310994 221656
rect 311102 221568 311282 221656
rect 311390 221568 311570 221656
rect 311678 221568 311858 221656
rect 311966 221568 312146 221656
rect 312254 221568 312434 221656
rect 312542 221568 312722 221656
rect 312830 221568 313010 221656
rect 325310 221568 325490 221656
rect 325598 221568 325778 221656
rect 325886 221568 326066 221656
rect 326174 221568 326354 221656
rect 326462 221568 326642 221656
rect 326750 221568 326930 221656
rect 327038 221568 327218 221656
rect 327326 221568 327506 221656
rect 339806 221568 339986 221656
rect 340094 221568 340274 221656
rect 340382 221568 340562 221656
rect 340670 221568 340850 221656
rect 340958 221568 341138 221656
rect 341246 221568 341426 221656
rect 341534 221568 341714 221656
rect 341822 221568 342002 221656
rect 354302 221568 354482 221656
rect 354590 221568 354770 221656
rect 354878 221568 355058 221656
rect 355166 221568 355346 221656
rect 355454 221568 355634 221656
rect 355742 221568 355922 221656
rect 356030 221568 356210 221656
rect 356318 221568 356498 221656
rect 368798 221568 368978 221656
rect 369086 221568 369266 221656
rect 369374 221568 369554 221656
rect 369662 221568 369842 221656
rect 369950 221568 370130 221656
rect 370238 221568 370418 221656
rect 370526 221568 370706 221656
rect 370814 221568 370994 221656
rect 383294 221568 383474 221656
rect 383582 221568 383762 221656
rect 383870 221568 384050 221656
rect 384158 221568 384338 221656
rect 384446 221568 384626 221656
rect 384734 221568 384914 221656
rect 385022 221568 385202 221656
rect 385310 221568 385490 221656
rect 397790 221568 397970 221656
rect 398078 221568 398258 221656
rect 398366 221568 398546 221656
rect 398654 221568 398834 221656
rect 398942 221568 399122 221656
rect 399230 221568 399410 221656
rect 399518 221568 399698 221656
rect 399806 221568 399986 221656
rect 412286 221568 412466 221656
rect 412574 221568 412754 221656
rect 412862 221568 413042 221656
rect 413150 221568 413330 221656
rect 413438 221568 413618 221656
rect 413726 221568 413906 221656
rect 414014 221568 414194 221656
rect 414302 221568 414482 221656
rect 426782 221568 426962 221656
rect 427070 221568 427250 221656
rect 427358 221568 427538 221656
rect 427646 221568 427826 221656
rect 427934 221568 428114 221656
rect 428222 221568 428402 221656
rect 428510 221568 428690 221656
rect 428798 221568 428978 221656
rect 441278 221568 441458 221656
rect 441566 221568 441746 221656
rect 441854 221568 442034 221656
rect 442142 221568 442322 221656
rect 442430 221568 442610 221656
rect 442718 221568 442898 221656
rect 443006 221568 443186 221656
rect 443294 221568 443474 221656
rect 455774 221568 455954 221656
rect 456062 221568 456242 221656
rect 456350 221568 456530 221656
rect 456638 221568 456818 221656
rect 456926 221568 457106 221656
rect 457214 221568 457394 221656
rect 457502 221568 457682 221656
rect 457790 221568 457970 221656
rect 180350 221352 180530 221440
rect 180638 221352 180818 221440
rect 180926 221352 181106 221440
rect 181214 221352 181394 221440
rect 181502 221352 181682 221440
rect 181790 221352 181970 221440
rect 182078 221352 182258 221440
rect 182366 221352 182546 221440
rect 194846 221352 195026 221440
rect 195134 221352 195314 221440
rect 195422 221352 195602 221440
rect 195710 221352 195890 221440
rect 195998 221352 196178 221440
rect 196286 221352 196466 221440
rect 196574 221352 196754 221440
rect 196862 221352 197042 221440
rect 209342 221352 209522 221440
rect 209630 221352 209810 221440
rect 209918 221352 210098 221440
rect 210206 221352 210386 221440
rect 210494 221352 210674 221440
rect 210782 221352 210962 221440
rect 211070 221352 211250 221440
rect 211358 221352 211538 221440
rect 223838 221352 224018 221440
rect 224126 221352 224306 221440
rect 224414 221352 224594 221440
rect 224702 221352 224882 221440
rect 224990 221352 225170 221440
rect 225278 221352 225458 221440
rect 225566 221352 225746 221440
rect 225854 221352 226034 221440
rect 238334 221352 238514 221440
rect 238622 221352 238802 221440
rect 238910 221352 239090 221440
rect 239198 221352 239378 221440
rect 239486 221352 239666 221440
rect 239774 221352 239954 221440
rect 240062 221352 240242 221440
rect 240350 221352 240530 221440
rect 252830 221352 253010 221440
rect 253118 221352 253298 221440
rect 253406 221352 253586 221440
rect 253694 221352 253874 221440
rect 253982 221352 254162 221440
rect 254270 221352 254450 221440
rect 254558 221352 254738 221440
rect 254846 221352 255026 221440
rect 267326 221352 267506 221440
rect 267614 221352 267794 221440
rect 267902 221352 268082 221440
rect 268190 221352 268370 221440
rect 268478 221352 268658 221440
rect 268766 221352 268946 221440
rect 269054 221352 269234 221440
rect 269342 221352 269522 221440
rect 281822 221352 282002 221440
rect 282110 221352 282290 221440
rect 282398 221352 282578 221440
rect 282686 221352 282866 221440
rect 282974 221352 283154 221440
rect 283262 221352 283442 221440
rect 283550 221352 283730 221440
rect 283838 221352 284018 221440
rect 296318 221352 296498 221440
rect 296606 221352 296786 221440
rect 296894 221352 297074 221440
rect 297182 221352 297362 221440
rect 297470 221352 297650 221440
rect 297758 221352 297938 221440
rect 298046 221352 298226 221440
rect 298334 221352 298514 221440
rect 310814 221352 310994 221440
rect 311102 221352 311282 221440
rect 311390 221352 311570 221440
rect 311678 221352 311858 221440
rect 311966 221352 312146 221440
rect 312254 221352 312434 221440
rect 312542 221352 312722 221440
rect 312830 221352 313010 221440
rect 325310 221352 325490 221440
rect 325598 221352 325778 221440
rect 325886 221352 326066 221440
rect 326174 221352 326354 221440
rect 326462 221352 326642 221440
rect 326750 221352 326930 221440
rect 327038 221352 327218 221440
rect 327326 221352 327506 221440
rect 339806 221352 339986 221440
rect 340094 221352 340274 221440
rect 340382 221352 340562 221440
rect 340670 221352 340850 221440
rect 340958 221352 341138 221440
rect 341246 221352 341426 221440
rect 341534 221352 341714 221440
rect 341822 221352 342002 221440
rect 354302 221352 354482 221440
rect 354590 221352 354770 221440
rect 354878 221352 355058 221440
rect 355166 221352 355346 221440
rect 355454 221352 355634 221440
rect 355742 221352 355922 221440
rect 356030 221352 356210 221440
rect 356318 221352 356498 221440
rect 368798 221352 368978 221440
rect 369086 221352 369266 221440
rect 369374 221352 369554 221440
rect 369662 221352 369842 221440
rect 369950 221352 370130 221440
rect 370238 221352 370418 221440
rect 370526 221352 370706 221440
rect 370814 221352 370994 221440
rect 383294 221352 383474 221440
rect 383582 221352 383762 221440
rect 383870 221352 384050 221440
rect 384158 221352 384338 221440
rect 384446 221352 384626 221440
rect 384734 221352 384914 221440
rect 385022 221352 385202 221440
rect 385310 221352 385490 221440
rect 397790 221352 397970 221440
rect 398078 221352 398258 221440
rect 398366 221352 398546 221440
rect 398654 221352 398834 221440
rect 398942 221352 399122 221440
rect 399230 221352 399410 221440
rect 399518 221352 399698 221440
rect 399806 221352 399986 221440
rect 412286 221352 412466 221440
rect 412574 221352 412754 221440
rect 412862 221352 413042 221440
rect 413150 221352 413330 221440
rect 413438 221352 413618 221440
rect 413726 221352 413906 221440
rect 414014 221352 414194 221440
rect 414302 221352 414482 221440
rect 426782 221352 426962 221440
rect 427070 221352 427250 221440
rect 427358 221352 427538 221440
rect 427646 221352 427826 221440
rect 427934 221352 428114 221440
rect 428222 221352 428402 221440
rect 428510 221352 428690 221440
rect 428798 221352 428978 221440
rect 441278 221352 441458 221440
rect 441566 221352 441746 221440
rect 441854 221352 442034 221440
rect 442142 221352 442322 221440
rect 442430 221352 442610 221440
rect 442718 221352 442898 221440
rect 443006 221352 443186 221440
rect 443294 221352 443474 221440
rect 455774 221352 455954 221440
rect 456062 221352 456242 221440
rect 456350 221352 456530 221440
rect 456638 221352 456818 221440
rect 456926 221352 457106 221440
rect 457214 221352 457394 221440
rect 457502 221352 457682 221440
rect 457790 221352 457970 221440
rect 180350 220876 180530 220964
rect 180638 220876 180818 220964
rect 180926 220876 181106 220964
rect 181214 220876 181394 220964
rect 181502 220876 181682 220964
rect 181790 220876 181970 220964
rect 182078 220876 182258 220964
rect 182366 220876 182546 220964
rect 194846 220876 195026 220964
rect 195134 220876 195314 220964
rect 195422 220876 195602 220964
rect 195710 220876 195890 220964
rect 195998 220876 196178 220964
rect 196286 220876 196466 220964
rect 196574 220876 196754 220964
rect 196862 220876 197042 220964
rect 209342 220876 209522 220964
rect 209630 220876 209810 220964
rect 209918 220876 210098 220964
rect 210206 220876 210386 220964
rect 210494 220876 210674 220964
rect 210782 220876 210962 220964
rect 211070 220876 211250 220964
rect 211358 220876 211538 220964
rect 223838 220876 224018 220964
rect 224126 220876 224306 220964
rect 224414 220876 224594 220964
rect 224702 220876 224882 220964
rect 224990 220876 225170 220964
rect 225278 220876 225458 220964
rect 225566 220876 225746 220964
rect 225854 220876 226034 220964
rect 238334 220876 238514 220964
rect 238622 220876 238802 220964
rect 238910 220876 239090 220964
rect 239198 220876 239378 220964
rect 239486 220876 239666 220964
rect 239774 220876 239954 220964
rect 240062 220876 240242 220964
rect 240350 220876 240530 220964
rect 252830 220876 253010 220964
rect 253118 220876 253298 220964
rect 253406 220876 253586 220964
rect 253694 220876 253874 220964
rect 253982 220876 254162 220964
rect 254270 220876 254450 220964
rect 254558 220876 254738 220964
rect 254846 220876 255026 220964
rect 267326 220876 267506 220964
rect 267614 220876 267794 220964
rect 267902 220876 268082 220964
rect 268190 220876 268370 220964
rect 268478 220876 268658 220964
rect 268766 220876 268946 220964
rect 269054 220876 269234 220964
rect 269342 220876 269522 220964
rect 281822 220876 282002 220964
rect 282110 220876 282290 220964
rect 282398 220876 282578 220964
rect 282686 220876 282866 220964
rect 282974 220876 283154 220964
rect 283262 220876 283442 220964
rect 283550 220876 283730 220964
rect 283838 220876 284018 220964
rect 296318 220876 296498 220964
rect 296606 220876 296786 220964
rect 296894 220876 297074 220964
rect 297182 220876 297362 220964
rect 297470 220876 297650 220964
rect 297758 220876 297938 220964
rect 298046 220876 298226 220964
rect 298334 220876 298514 220964
rect 310814 220876 310994 220964
rect 311102 220876 311282 220964
rect 311390 220876 311570 220964
rect 311678 220876 311858 220964
rect 311966 220876 312146 220964
rect 312254 220876 312434 220964
rect 312542 220876 312722 220964
rect 312830 220876 313010 220964
rect 325310 220876 325490 220964
rect 325598 220876 325778 220964
rect 325886 220876 326066 220964
rect 326174 220876 326354 220964
rect 326462 220876 326642 220964
rect 326750 220876 326930 220964
rect 327038 220876 327218 220964
rect 327326 220876 327506 220964
rect 339806 220876 339986 220964
rect 340094 220876 340274 220964
rect 340382 220876 340562 220964
rect 340670 220876 340850 220964
rect 340958 220876 341138 220964
rect 341246 220876 341426 220964
rect 341534 220876 341714 220964
rect 341822 220876 342002 220964
rect 354302 220876 354482 220964
rect 354590 220876 354770 220964
rect 354878 220876 355058 220964
rect 355166 220876 355346 220964
rect 355454 220876 355634 220964
rect 355742 220876 355922 220964
rect 356030 220876 356210 220964
rect 356318 220876 356498 220964
rect 368798 220876 368978 220964
rect 369086 220876 369266 220964
rect 369374 220876 369554 220964
rect 369662 220876 369842 220964
rect 369950 220876 370130 220964
rect 370238 220876 370418 220964
rect 370526 220876 370706 220964
rect 370814 220876 370994 220964
rect 383294 220876 383474 220964
rect 383582 220876 383762 220964
rect 383870 220876 384050 220964
rect 384158 220876 384338 220964
rect 384446 220876 384626 220964
rect 384734 220876 384914 220964
rect 385022 220876 385202 220964
rect 385310 220876 385490 220964
rect 397790 220876 397970 220964
rect 398078 220876 398258 220964
rect 398366 220876 398546 220964
rect 398654 220876 398834 220964
rect 398942 220876 399122 220964
rect 399230 220876 399410 220964
rect 399518 220876 399698 220964
rect 399806 220876 399986 220964
rect 412286 220876 412466 220964
rect 412574 220876 412754 220964
rect 412862 220876 413042 220964
rect 413150 220876 413330 220964
rect 413438 220876 413618 220964
rect 413726 220876 413906 220964
rect 414014 220876 414194 220964
rect 414302 220876 414482 220964
rect 426782 220876 426962 220964
rect 427070 220876 427250 220964
rect 427358 220876 427538 220964
rect 427646 220876 427826 220964
rect 427934 220876 428114 220964
rect 428222 220876 428402 220964
rect 428510 220876 428690 220964
rect 428798 220876 428978 220964
rect 441278 220876 441458 220964
rect 441566 220876 441746 220964
rect 441854 220876 442034 220964
rect 442142 220876 442322 220964
rect 442430 220876 442610 220964
rect 442718 220876 442898 220964
rect 443006 220876 443186 220964
rect 443294 220876 443474 220964
rect 455774 220876 455954 220964
rect 456062 220876 456242 220964
rect 456350 220876 456530 220964
rect 456638 220876 456818 220964
rect 456926 220876 457106 220964
rect 457214 220876 457394 220964
rect 457502 220876 457682 220964
rect 457790 220876 457970 220964
rect 180350 220660 180530 220748
rect 180638 220660 180818 220748
rect 180926 220660 181106 220748
rect 181214 220660 181394 220748
rect 181502 220660 181682 220748
rect 181790 220660 181970 220748
rect 182078 220660 182258 220748
rect 182366 220660 182546 220748
rect 194846 220660 195026 220748
rect 195134 220660 195314 220748
rect 195422 220660 195602 220748
rect 195710 220660 195890 220748
rect 195998 220660 196178 220748
rect 196286 220660 196466 220748
rect 196574 220660 196754 220748
rect 196862 220660 197042 220748
rect 209342 220660 209522 220748
rect 209630 220660 209810 220748
rect 209918 220660 210098 220748
rect 210206 220660 210386 220748
rect 210494 220660 210674 220748
rect 210782 220660 210962 220748
rect 211070 220660 211250 220748
rect 211358 220660 211538 220748
rect 223838 220660 224018 220748
rect 224126 220660 224306 220748
rect 224414 220660 224594 220748
rect 224702 220660 224882 220748
rect 224990 220660 225170 220748
rect 225278 220660 225458 220748
rect 225566 220660 225746 220748
rect 225854 220660 226034 220748
rect 238334 220660 238514 220748
rect 238622 220660 238802 220748
rect 238910 220660 239090 220748
rect 239198 220660 239378 220748
rect 239486 220660 239666 220748
rect 239774 220660 239954 220748
rect 240062 220660 240242 220748
rect 240350 220660 240530 220748
rect 252830 220660 253010 220748
rect 253118 220660 253298 220748
rect 253406 220660 253586 220748
rect 253694 220660 253874 220748
rect 253982 220660 254162 220748
rect 254270 220660 254450 220748
rect 254558 220660 254738 220748
rect 254846 220660 255026 220748
rect 267326 220660 267506 220748
rect 267614 220660 267794 220748
rect 267902 220660 268082 220748
rect 268190 220660 268370 220748
rect 268478 220660 268658 220748
rect 268766 220660 268946 220748
rect 269054 220660 269234 220748
rect 269342 220660 269522 220748
rect 281822 220660 282002 220748
rect 282110 220660 282290 220748
rect 282398 220660 282578 220748
rect 282686 220660 282866 220748
rect 282974 220660 283154 220748
rect 283262 220660 283442 220748
rect 283550 220660 283730 220748
rect 283838 220660 284018 220748
rect 296318 220660 296498 220748
rect 296606 220660 296786 220748
rect 296894 220660 297074 220748
rect 297182 220660 297362 220748
rect 297470 220660 297650 220748
rect 297758 220660 297938 220748
rect 298046 220660 298226 220748
rect 298334 220660 298514 220748
rect 310814 220660 310994 220748
rect 311102 220660 311282 220748
rect 311390 220660 311570 220748
rect 311678 220660 311858 220748
rect 311966 220660 312146 220748
rect 312254 220660 312434 220748
rect 312542 220660 312722 220748
rect 312830 220660 313010 220748
rect 325310 220660 325490 220748
rect 325598 220660 325778 220748
rect 325886 220660 326066 220748
rect 326174 220660 326354 220748
rect 326462 220660 326642 220748
rect 326750 220660 326930 220748
rect 327038 220660 327218 220748
rect 327326 220660 327506 220748
rect 339806 220660 339986 220748
rect 340094 220660 340274 220748
rect 340382 220660 340562 220748
rect 340670 220660 340850 220748
rect 340958 220660 341138 220748
rect 341246 220660 341426 220748
rect 341534 220660 341714 220748
rect 341822 220660 342002 220748
rect 354302 220660 354482 220748
rect 354590 220660 354770 220748
rect 354878 220660 355058 220748
rect 355166 220660 355346 220748
rect 355454 220660 355634 220748
rect 355742 220660 355922 220748
rect 356030 220660 356210 220748
rect 356318 220660 356498 220748
rect 368798 220660 368978 220748
rect 369086 220660 369266 220748
rect 369374 220660 369554 220748
rect 369662 220660 369842 220748
rect 369950 220660 370130 220748
rect 370238 220660 370418 220748
rect 370526 220660 370706 220748
rect 370814 220660 370994 220748
rect 383294 220660 383474 220748
rect 383582 220660 383762 220748
rect 383870 220660 384050 220748
rect 384158 220660 384338 220748
rect 384446 220660 384626 220748
rect 384734 220660 384914 220748
rect 385022 220660 385202 220748
rect 385310 220660 385490 220748
rect 397790 220660 397970 220748
rect 398078 220660 398258 220748
rect 398366 220660 398546 220748
rect 398654 220660 398834 220748
rect 398942 220660 399122 220748
rect 399230 220660 399410 220748
rect 399518 220660 399698 220748
rect 399806 220660 399986 220748
rect 412286 220660 412466 220748
rect 412574 220660 412754 220748
rect 412862 220660 413042 220748
rect 413150 220660 413330 220748
rect 413438 220660 413618 220748
rect 413726 220660 413906 220748
rect 414014 220660 414194 220748
rect 414302 220660 414482 220748
rect 426782 220660 426962 220748
rect 427070 220660 427250 220748
rect 427358 220660 427538 220748
rect 427646 220660 427826 220748
rect 427934 220660 428114 220748
rect 428222 220660 428402 220748
rect 428510 220660 428690 220748
rect 428798 220660 428978 220748
rect 441278 220660 441458 220748
rect 441566 220660 441746 220748
rect 441854 220660 442034 220748
rect 442142 220660 442322 220748
rect 442430 220660 442610 220748
rect 442718 220660 442898 220748
rect 443006 220660 443186 220748
rect 443294 220660 443474 220748
rect 455774 220660 455954 220748
rect 456062 220660 456242 220748
rect 456350 220660 456530 220748
rect 456638 220660 456818 220748
rect 456926 220660 457106 220748
rect 457214 220660 457394 220748
rect 457502 220660 457682 220748
rect 457790 220660 457970 220748
rect 180350 206508 180530 206596
rect 180638 206508 180818 206596
rect 180926 206508 181106 206596
rect 181214 206508 181394 206596
rect 181502 206508 181682 206596
rect 181790 206508 181970 206596
rect 182078 206508 182258 206596
rect 182366 206508 182546 206596
rect 194846 206508 195026 206596
rect 195134 206508 195314 206596
rect 195422 206508 195602 206596
rect 195710 206508 195890 206596
rect 195998 206508 196178 206596
rect 196286 206508 196466 206596
rect 196574 206508 196754 206596
rect 196862 206508 197042 206596
rect 209342 206508 209522 206596
rect 209630 206508 209810 206596
rect 209918 206508 210098 206596
rect 210206 206508 210386 206596
rect 210494 206508 210674 206596
rect 210782 206508 210962 206596
rect 211070 206508 211250 206596
rect 211358 206508 211538 206596
rect 223838 206508 224018 206596
rect 224126 206508 224306 206596
rect 224414 206508 224594 206596
rect 224702 206508 224882 206596
rect 224990 206508 225170 206596
rect 225278 206508 225458 206596
rect 225566 206508 225746 206596
rect 225854 206508 226034 206596
rect 238334 206508 238514 206596
rect 238622 206508 238802 206596
rect 238910 206508 239090 206596
rect 239198 206508 239378 206596
rect 239486 206508 239666 206596
rect 239774 206508 239954 206596
rect 240062 206508 240242 206596
rect 240350 206508 240530 206596
rect 252830 206508 253010 206596
rect 253118 206508 253298 206596
rect 253406 206508 253586 206596
rect 253694 206508 253874 206596
rect 253982 206508 254162 206596
rect 254270 206508 254450 206596
rect 254558 206508 254738 206596
rect 254846 206508 255026 206596
rect 267326 206508 267506 206596
rect 267614 206508 267794 206596
rect 267902 206508 268082 206596
rect 268190 206508 268370 206596
rect 268478 206508 268658 206596
rect 268766 206508 268946 206596
rect 269054 206508 269234 206596
rect 269342 206508 269522 206596
rect 281822 206508 282002 206596
rect 282110 206508 282290 206596
rect 282398 206508 282578 206596
rect 282686 206508 282866 206596
rect 282974 206508 283154 206596
rect 283262 206508 283442 206596
rect 283550 206508 283730 206596
rect 283838 206508 284018 206596
rect 296318 206508 296498 206596
rect 296606 206508 296786 206596
rect 296894 206508 297074 206596
rect 297182 206508 297362 206596
rect 297470 206508 297650 206596
rect 297758 206508 297938 206596
rect 298046 206508 298226 206596
rect 298334 206508 298514 206596
rect 310814 206508 310994 206596
rect 311102 206508 311282 206596
rect 311390 206508 311570 206596
rect 311678 206508 311858 206596
rect 311966 206508 312146 206596
rect 312254 206508 312434 206596
rect 312542 206508 312722 206596
rect 312830 206508 313010 206596
rect 325310 206508 325490 206596
rect 325598 206508 325778 206596
rect 325886 206508 326066 206596
rect 326174 206508 326354 206596
rect 326462 206508 326642 206596
rect 326750 206508 326930 206596
rect 327038 206508 327218 206596
rect 327326 206508 327506 206596
rect 339806 206508 339986 206596
rect 340094 206508 340274 206596
rect 340382 206508 340562 206596
rect 340670 206508 340850 206596
rect 340958 206508 341138 206596
rect 341246 206508 341426 206596
rect 341534 206508 341714 206596
rect 341822 206508 342002 206596
rect 354302 206508 354482 206596
rect 354590 206508 354770 206596
rect 354878 206508 355058 206596
rect 355166 206508 355346 206596
rect 355454 206508 355634 206596
rect 355742 206508 355922 206596
rect 356030 206508 356210 206596
rect 356318 206508 356498 206596
rect 368798 206508 368978 206596
rect 369086 206508 369266 206596
rect 369374 206508 369554 206596
rect 369662 206508 369842 206596
rect 369950 206508 370130 206596
rect 370238 206508 370418 206596
rect 370526 206508 370706 206596
rect 370814 206508 370994 206596
rect 383294 206508 383474 206596
rect 383582 206508 383762 206596
rect 383870 206508 384050 206596
rect 384158 206508 384338 206596
rect 384446 206508 384626 206596
rect 384734 206508 384914 206596
rect 385022 206508 385202 206596
rect 385310 206508 385490 206596
rect 397790 206508 397970 206596
rect 398078 206508 398258 206596
rect 398366 206508 398546 206596
rect 398654 206508 398834 206596
rect 398942 206508 399122 206596
rect 399230 206508 399410 206596
rect 399518 206508 399698 206596
rect 399806 206508 399986 206596
rect 412286 206508 412466 206596
rect 412574 206508 412754 206596
rect 412862 206508 413042 206596
rect 413150 206508 413330 206596
rect 413438 206508 413618 206596
rect 413726 206508 413906 206596
rect 414014 206508 414194 206596
rect 414302 206508 414482 206596
rect 426782 206508 426962 206596
rect 427070 206508 427250 206596
rect 427358 206508 427538 206596
rect 427646 206508 427826 206596
rect 427934 206508 428114 206596
rect 428222 206508 428402 206596
rect 428510 206508 428690 206596
rect 428798 206508 428978 206596
rect 441278 206508 441458 206596
rect 441566 206508 441746 206596
rect 441854 206508 442034 206596
rect 442142 206508 442322 206596
rect 442430 206508 442610 206596
rect 442718 206508 442898 206596
rect 443006 206508 443186 206596
rect 443294 206508 443474 206596
rect 455774 206508 455954 206596
rect 456062 206508 456242 206596
rect 456350 206508 456530 206596
rect 456638 206508 456818 206596
rect 456926 206508 457106 206596
rect 457214 206508 457394 206596
rect 457502 206508 457682 206596
rect 457790 206508 457970 206596
rect 180350 206292 180530 206380
rect 180638 206292 180818 206380
rect 180926 206292 181106 206380
rect 181214 206292 181394 206380
rect 181502 206292 181682 206380
rect 181790 206292 181970 206380
rect 182078 206292 182258 206380
rect 182366 206292 182546 206380
rect 194846 206292 195026 206380
rect 195134 206292 195314 206380
rect 195422 206292 195602 206380
rect 195710 206292 195890 206380
rect 195998 206292 196178 206380
rect 196286 206292 196466 206380
rect 196574 206292 196754 206380
rect 196862 206292 197042 206380
rect 209342 206292 209522 206380
rect 209630 206292 209810 206380
rect 209918 206292 210098 206380
rect 210206 206292 210386 206380
rect 210494 206292 210674 206380
rect 210782 206292 210962 206380
rect 211070 206292 211250 206380
rect 211358 206292 211538 206380
rect 223838 206292 224018 206380
rect 224126 206292 224306 206380
rect 224414 206292 224594 206380
rect 224702 206292 224882 206380
rect 224990 206292 225170 206380
rect 225278 206292 225458 206380
rect 225566 206292 225746 206380
rect 225854 206292 226034 206380
rect 238334 206292 238514 206380
rect 238622 206292 238802 206380
rect 238910 206292 239090 206380
rect 239198 206292 239378 206380
rect 239486 206292 239666 206380
rect 239774 206292 239954 206380
rect 240062 206292 240242 206380
rect 240350 206292 240530 206380
rect 252830 206292 253010 206380
rect 253118 206292 253298 206380
rect 253406 206292 253586 206380
rect 253694 206292 253874 206380
rect 253982 206292 254162 206380
rect 254270 206292 254450 206380
rect 254558 206292 254738 206380
rect 254846 206292 255026 206380
rect 267326 206292 267506 206380
rect 267614 206292 267794 206380
rect 267902 206292 268082 206380
rect 268190 206292 268370 206380
rect 268478 206292 268658 206380
rect 268766 206292 268946 206380
rect 269054 206292 269234 206380
rect 269342 206292 269522 206380
rect 281822 206292 282002 206380
rect 282110 206292 282290 206380
rect 282398 206292 282578 206380
rect 282686 206292 282866 206380
rect 282974 206292 283154 206380
rect 283262 206292 283442 206380
rect 283550 206292 283730 206380
rect 283838 206292 284018 206380
rect 296318 206292 296498 206380
rect 296606 206292 296786 206380
rect 296894 206292 297074 206380
rect 297182 206292 297362 206380
rect 297470 206292 297650 206380
rect 297758 206292 297938 206380
rect 298046 206292 298226 206380
rect 298334 206292 298514 206380
rect 310814 206292 310994 206380
rect 311102 206292 311282 206380
rect 311390 206292 311570 206380
rect 311678 206292 311858 206380
rect 311966 206292 312146 206380
rect 312254 206292 312434 206380
rect 312542 206292 312722 206380
rect 312830 206292 313010 206380
rect 325310 206292 325490 206380
rect 325598 206292 325778 206380
rect 325886 206292 326066 206380
rect 326174 206292 326354 206380
rect 326462 206292 326642 206380
rect 326750 206292 326930 206380
rect 327038 206292 327218 206380
rect 327326 206292 327506 206380
rect 339806 206292 339986 206380
rect 340094 206292 340274 206380
rect 340382 206292 340562 206380
rect 340670 206292 340850 206380
rect 340958 206292 341138 206380
rect 341246 206292 341426 206380
rect 341534 206292 341714 206380
rect 341822 206292 342002 206380
rect 354302 206292 354482 206380
rect 354590 206292 354770 206380
rect 354878 206292 355058 206380
rect 355166 206292 355346 206380
rect 355454 206292 355634 206380
rect 355742 206292 355922 206380
rect 356030 206292 356210 206380
rect 356318 206292 356498 206380
rect 368798 206292 368978 206380
rect 369086 206292 369266 206380
rect 369374 206292 369554 206380
rect 369662 206292 369842 206380
rect 369950 206292 370130 206380
rect 370238 206292 370418 206380
rect 370526 206292 370706 206380
rect 370814 206292 370994 206380
rect 383294 206292 383474 206380
rect 383582 206292 383762 206380
rect 383870 206292 384050 206380
rect 384158 206292 384338 206380
rect 384446 206292 384626 206380
rect 384734 206292 384914 206380
rect 385022 206292 385202 206380
rect 385310 206292 385490 206380
rect 397790 206292 397970 206380
rect 398078 206292 398258 206380
rect 398366 206292 398546 206380
rect 398654 206292 398834 206380
rect 398942 206292 399122 206380
rect 399230 206292 399410 206380
rect 399518 206292 399698 206380
rect 399806 206292 399986 206380
rect 412286 206292 412466 206380
rect 412574 206292 412754 206380
rect 412862 206292 413042 206380
rect 413150 206292 413330 206380
rect 413438 206292 413618 206380
rect 413726 206292 413906 206380
rect 414014 206292 414194 206380
rect 414302 206292 414482 206380
rect 426782 206292 426962 206380
rect 427070 206292 427250 206380
rect 427358 206292 427538 206380
rect 427646 206292 427826 206380
rect 427934 206292 428114 206380
rect 428222 206292 428402 206380
rect 428510 206292 428690 206380
rect 428798 206292 428978 206380
rect 441278 206292 441458 206380
rect 441566 206292 441746 206380
rect 441854 206292 442034 206380
rect 442142 206292 442322 206380
rect 442430 206292 442610 206380
rect 442718 206292 442898 206380
rect 443006 206292 443186 206380
rect 443294 206292 443474 206380
rect 455774 206292 455954 206380
rect 456062 206292 456242 206380
rect 456350 206292 456530 206380
rect 456638 206292 456818 206380
rect 456926 206292 457106 206380
rect 457214 206292 457394 206380
rect 457502 206292 457682 206380
rect 457790 206292 457970 206380
rect 180350 205816 180530 205904
rect 180638 205816 180818 205904
rect 180926 205816 181106 205904
rect 181214 205816 181394 205904
rect 181502 205816 181682 205904
rect 181790 205816 181970 205904
rect 182078 205816 182258 205904
rect 182366 205816 182546 205904
rect 194846 205816 195026 205904
rect 195134 205816 195314 205904
rect 195422 205816 195602 205904
rect 195710 205816 195890 205904
rect 195998 205816 196178 205904
rect 196286 205816 196466 205904
rect 196574 205816 196754 205904
rect 196862 205816 197042 205904
rect 209342 205816 209522 205904
rect 209630 205816 209810 205904
rect 209918 205816 210098 205904
rect 210206 205816 210386 205904
rect 210494 205816 210674 205904
rect 210782 205816 210962 205904
rect 211070 205816 211250 205904
rect 211358 205816 211538 205904
rect 223838 205816 224018 205904
rect 224126 205816 224306 205904
rect 224414 205816 224594 205904
rect 224702 205816 224882 205904
rect 224990 205816 225170 205904
rect 225278 205816 225458 205904
rect 225566 205816 225746 205904
rect 225854 205816 226034 205904
rect 238334 205816 238514 205904
rect 238622 205816 238802 205904
rect 238910 205816 239090 205904
rect 239198 205816 239378 205904
rect 239486 205816 239666 205904
rect 239774 205816 239954 205904
rect 240062 205816 240242 205904
rect 240350 205816 240530 205904
rect 252830 205816 253010 205904
rect 253118 205816 253298 205904
rect 253406 205816 253586 205904
rect 253694 205816 253874 205904
rect 253982 205816 254162 205904
rect 254270 205816 254450 205904
rect 254558 205816 254738 205904
rect 254846 205816 255026 205904
rect 267326 205816 267506 205904
rect 267614 205816 267794 205904
rect 267902 205816 268082 205904
rect 268190 205816 268370 205904
rect 268478 205816 268658 205904
rect 268766 205816 268946 205904
rect 269054 205816 269234 205904
rect 269342 205816 269522 205904
rect 281822 205816 282002 205904
rect 282110 205816 282290 205904
rect 282398 205816 282578 205904
rect 282686 205816 282866 205904
rect 282974 205816 283154 205904
rect 283262 205816 283442 205904
rect 283550 205816 283730 205904
rect 283838 205816 284018 205904
rect 296318 205816 296498 205904
rect 296606 205816 296786 205904
rect 296894 205816 297074 205904
rect 297182 205816 297362 205904
rect 297470 205816 297650 205904
rect 297758 205816 297938 205904
rect 298046 205816 298226 205904
rect 298334 205816 298514 205904
rect 310814 205816 310994 205904
rect 311102 205816 311282 205904
rect 311390 205816 311570 205904
rect 311678 205816 311858 205904
rect 311966 205816 312146 205904
rect 312254 205816 312434 205904
rect 312542 205816 312722 205904
rect 312830 205816 313010 205904
rect 325310 205816 325490 205904
rect 325598 205816 325778 205904
rect 325886 205816 326066 205904
rect 326174 205816 326354 205904
rect 326462 205816 326642 205904
rect 326750 205816 326930 205904
rect 327038 205816 327218 205904
rect 327326 205816 327506 205904
rect 339806 205816 339986 205904
rect 340094 205816 340274 205904
rect 340382 205816 340562 205904
rect 340670 205816 340850 205904
rect 340958 205816 341138 205904
rect 341246 205816 341426 205904
rect 341534 205816 341714 205904
rect 341822 205816 342002 205904
rect 354302 205816 354482 205904
rect 354590 205816 354770 205904
rect 354878 205816 355058 205904
rect 355166 205816 355346 205904
rect 355454 205816 355634 205904
rect 355742 205816 355922 205904
rect 356030 205816 356210 205904
rect 356318 205816 356498 205904
rect 368798 205816 368978 205904
rect 369086 205816 369266 205904
rect 369374 205816 369554 205904
rect 369662 205816 369842 205904
rect 369950 205816 370130 205904
rect 370238 205816 370418 205904
rect 370526 205816 370706 205904
rect 370814 205816 370994 205904
rect 383294 205816 383474 205904
rect 383582 205816 383762 205904
rect 383870 205816 384050 205904
rect 384158 205816 384338 205904
rect 384446 205816 384626 205904
rect 384734 205816 384914 205904
rect 385022 205816 385202 205904
rect 385310 205816 385490 205904
rect 397790 205816 397970 205904
rect 398078 205816 398258 205904
rect 398366 205816 398546 205904
rect 398654 205816 398834 205904
rect 398942 205816 399122 205904
rect 399230 205816 399410 205904
rect 399518 205816 399698 205904
rect 399806 205816 399986 205904
rect 412286 205816 412466 205904
rect 412574 205816 412754 205904
rect 412862 205816 413042 205904
rect 413150 205816 413330 205904
rect 413438 205816 413618 205904
rect 413726 205816 413906 205904
rect 414014 205816 414194 205904
rect 414302 205816 414482 205904
rect 426782 205816 426962 205904
rect 427070 205816 427250 205904
rect 427358 205816 427538 205904
rect 427646 205816 427826 205904
rect 427934 205816 428114 205904
rect 428222 205816 428402 205904
rect 428510 205816 428690 205904
rect 428798 205816 428978 205904
rect 441278 205816 441458 205904
rect 441566 205816 441746 205904
rect 441854 205816 442034 205904
rect 442142 205816 442322 205904
rect 442430 205816 442610 205904
rect 442718 205816 442898 205904
rect 443006 205816 443186 205904
rect 443294 205816 443474 205904
rect 455774 205816 455954 205904
rect 456062 205816 456242 205904
rect 456350 205816 456530 205904
rect 456638 205816 456818 205904
rect 456926 205816 457106 205904
rect 457214 205816 457394 205904
rect 457502 205816 457682 205904
rect 457790 205816 457970 205904
rect 180350 205600 180530 205688
rect 180638 205600 180818 205688
rect 180926 205600 181106 205688
rect 181214 205600 181394 205688
rect 181502 205600 181682 205688
rect 181790 205600 181970 205688
rect 182078 205600 182258 205688
rect 182366 205600 182546 205688
rect 194846 205600 195026 205688
rect 195134 205600 195314 205688
rect 195422 205600 195602 205688
rect 195710 205600 195890 205688
rect 195998 205600 196178 205688
rect 196286 205600 196466 205688
rect 196574 205600 196754 205688
rect 196862 205600 197042 205688
rect 209342 205600 209522 205688
rect 209630 205600 209810 205688
rect 209918 205600 210098 205688
rect 210206 205600 210386 205688
rect 210494 205600 210674 205688
rect 210782 205600 210962 205688
rect 211070 205600 211250 205688
rect 211358 205600 211538 205688
rect 223838 205600 224018 205688
rect 224126 205600 224306 205688
rect 224414 205600 224594 205688
rect 224702 205600 224882 205688
rect 224990 205600 225170 205688
rect 225278 205600 225458 205688
rect 225566 205600 225746 205688
rect 225854 205600 226034 205688
rect 238334 205600 238514 205688
rect 238622 205600 238802 205688
rect 238910 205600 239090 205688
rect 239198 205600 239378 205688
rect 239486 205600 239666 205688
rect 239774 205600 239954 205688
rect 240062 205600 240242 205688
rect 240350 205600 240530 205688
rect 252830 205600 253010 205688
rect 253118 205600 253298 205688
rect 253406 205600 253586 205688
rect 253694 205600 253874 205688
rect 253982 205600 254162 205688
rect 254270 205600 254450 205688
rect 254558 205600 254738 205688
rect 254846 205600 255026 205688
rect 267326 205600 267506 205688
rect 267614 205600 267794 205688
rect 267902 205600 268082 205688
rect 268190 205600 268370 205688
rect 268478 205600 268658 205688
rect 268766 205600 268946 205688
rect 269054 205600 269234 205688
rect 269342 205600 269522 205688
rect 281822 205600 282002 205688
rect 282110 205600 282290 205688
rect 282398 205600 282578 205688
rect 282686 205600 282866 205688
rect 282974 205600 283154 205688
rect 283262 205600 283442 205688
rect 283550 205600 283730 205688
rect 283838 205600 284018 205688
rect 296318 205600 296498 205688
rect 296606 205600 296786 205688
rect 296894 205600 297074 205688
rect 297182 205600 297362 205688
rect 297470 205600 297650 205688
rect 297758 205600 297938 205688
rect 298046 205600 298226 205688
rect 298334 205600 298514 205688
rect 310814 205600 310994 205688
rect 311102 205600 311282 205688
rect 311390 205600 311570 205688
rect 311678 205600 311858 205688
rect 311966 205600 312146 205688
rect 312254 205600 312434 205688
rect 312542 205600 312722 205688
rect 312830 205600 313010 205688
rect 325310 205600 325490 205688
rect 325598 205600 325778 205688
rect 325886 205600 326066 205688
rect 326174 205600 326354 205688
rect 326462 205600 326642 205688
rect 326750 205600 326930 205688
rect 327038 205600 327218 205688
rect 327326 205600 327506 205688
rect 339806 205600 339986 205688
rect 340094 205600 340274 205688
rect 340382 205600 340562 205688
rect 340670 205600 340850 205688
rect 340958 205600 341138 205688
rect 341246 205600 341426 205688
rect 341534 205600 341714 205688
rect 341822 205600 342002 205688
rect 354302 205600 354482 205688
rect 354590 205600 354770 205688
rect 354878 205600 355058 205688
rect 355166 205600 355346 205688
rect 355454 205600 355634 205688
rect 355742 205600 355922 205688
rect 356030 205600 356210 205688
rect 356318 205600 356498 205688
rect 368798 205600 368978 205688
rect 369086 205600 369266 205688
rect 369374 205600 369554 205688
rect 369662 205600 369842 205688
rect 369950 205600 370130 205688
rect 370238 205600 370418 205688
rect 370526 205600 370706 205688
rect 370814 205600 370994 205688
rect 383294 205600 383474 205688
rect 383582 205600 383762 205688
rect 383870 205600 384050 205688
rect 384158 205600 384338 205688
rect 384446 205600 384626 205688
rect 384734 205600 384914 205688
rect 385022 205600 385202 205688
rect 385310 205600 385490 205688
rect 397790 205600 397970 205688
rect 398078 205600 398258 205688
rect 398366 205600 398546 205688
rect 398654 205600 398834 205688
rect 398942 205600 399122 205688
rect 399230 205600 399410 205688
rect 399518 205600 399698 205688
rect 399806 205600 399986 205688
rect 412286 205600 412466 205688
rect 412574 205600 412754 205688
rect 412862 205600 413042 205688
rect 413150 205600 413330 205688
rect 413438 205600 413618 205688
rect 413726 205600 413906 205688
rect 414014 205600 414194 205688
rect 414302 205600 414482 205688
rect 426782 205600 426962 205688
rect 427070 205600 427250 205688
rect 427358 205600 427538 205688
rect 427646 205600 427826 205688
rect 427934 205600 428114 205688
rect 428222 205600 428402 205688
rect 428510 205600 428690 205688
rect 428798 205600 428978 205688
rect 441278 205600 441458 205688
rect 441566 205600 441746 205688
rect 441854 205600 442034 205688
rect 442142 205600 442322 205688
rect 442430 205600 442610 205688
rect 442718 205600 442898 205688
rect 443006 205600 443186 205688
rect 443294 205600 443474 205688
rect 455774 205600 455954 205688
rect 456062 205600 456242 205688
rect 456350 205600 456530 205688
rect 456638 205600 456818 205688
rect 456926 205600 457106 205688
rect 457214 205600 457394 205688
rect 457502 205600 457682 205688
rect 457790 205600 457970 205688
rect 180350 191448 180530 191536
rect 180638 191448 180818 191536
rect 180926 191448 181106 191536
rect 181214 191448 181394 191536
rect 181502 191448 181682 191536
rect 181790 191448 181970 191536
rect 182078 191448 182258 191536
rect 182366 191448 182546 191536
rect 194846 191448 195026 191536
rect 195134 191448 195314 191536
rect 195422 191448 195602 191536
rect 195710 191448 195890 191536
rect 195998 191448 196178 191536
rect 196286 191448 196466 191536
rect 196574 191448 196754 191536
rect 196862 191448 197042 191536
rect 209342 191448 209522 191536
rect 209630 191448 209810 191536
rect 209918 191448 210098 191536
rect 210206 191448 210386 191536
rect 210494 191448 210674 191536
rect 210782 191448 210962 191536
rect 211070 191448 211250 191536
rect 211358 191448 211538 191536
rect 223838 191448 224018 191536
rect 224126 191448 224306 191536
rect 224414 191448 224594 191536
rect 224702 191448 224882 191536
rect 224990 191448 225170 191536
rect 225278 191448 225458 191536
rect 225566 191448 225746 191536
rect 225854 191448 226034 191536
rect 238334 191448 238514 191536
rect 238622 191448 238802 191536
rect 238910 191448 239090 191536
rect 239198 191448 239378 191536
rect 239486 191448 239666 191536
rect 239774 191448 239954 191536
rect 240062 191448 240242 191536
rect 240350 191448 240530 191536
rect 252830 191448 253010 191536
rect 253118 191448 253298 191536
rect 253406 191448 253586 191536
rect 253694 191448 253874 191536
rect 253982 191448 254162 191536
rect 254270 191448 254450 191536
rect 254558 191448 254738 191536
rect 254846 191448 255026 191536
rect 267326 191448 267506 191536
rect 267614 191448 267794 191536
rect 267902 191448 268082 191536
rect 268190 191448 268370 191536
rect 268478 191448 268658 191536
rect 268766 191448 268946 191536
rect 269054 191448 269234 191536
rect 269342 191448 269522 191536
rect 281822 191448 282002 191536
rect 282110 191448 282290 191536
rect 282398 191448 282578 191536
rect 282686 191448 282866 191536
rect 282974 191448 283154 191536
rect 283262 191448 283442 191536
rect 283550 191448 283730 191536
rect 283838 191448 284018 191536
rect 296318 191448 296498 191536
rect 296606 191448 296786 191536
rect 296894 191448 297074 191536
rect 297182 191448 297362 191536
rect 297470 191448 297650 191536
rect 297758 191448 297938 191536
rect 298046 191448 298226 191536
rect 298334 191448 298514 191536
rect 310814 191448 310994 191536
rect 311102 191448 311282 191536
rect 311390 191448 311570 191536
rect 311678 191448 311858 191536
rect 311966 191448 312146 191536
rect 312254 191448 312434 191536
rect 312542 191448 312722 191536
rect 312830 191448 313010 191536
rect 325310 191448 325490 191536
rect 325598 191448 325778 191536
rect 325886 191448 326066 191536
rect 326174 191448 326354 191536
rect 326462 191448 326642 191536
rect 326750 191448 326930 191536
rect 327038 191448 327218 191536
rect 327326 191448 327506 191536
rect 339806 191448 339986 191536
rect 340094 191448 340274 191536
rect 340382 191448 340562 191536
rect 340670 191448 340850 191536
rect 340958 191448 341138 191536
rect 341246 191448 341426 191536
rect 341534 191448 341714 191536
rect 341822 191448 342002 191536
rect 354302 191448 354482 191536
rect 354590 191448 354770 191536
rect 354878 191448 355058 191536
rect 355166 191448 355346 191536
rect 355454 191448 355634 191536
rect 355742 191448 355922 191536
rect 356030 191448 356210 191536
rect 356318 191448 356498 191536
rect 368798 191448 368978 191536
rect 369086 191448 369266 191536
rect 369374 191448 369554 191536
rect 369662 191448 369842 191536
rect 369950 191448 370130 191536
rect 370238 191448 370418 191536
rect 370526 191448 370706 191536
rect 370814 191448 370994 191536
rect 383294 191448 383474 191536
rect 383582 191448 383762 191536
rect 383870 191448 384050 191536
rect 384158 191448 384338 191536
rect 384446 191448 384626 191536
rect 384734 191448 384914 191536
rect 385022 191448 385202 191536
rect 385310 191448 385490 191536
rect 397790 191448 397970 191536
rect 398078 191448 398258 191536
rect 398366 191448 398546 191536
rect 398654 191448 398834 191536
rect 398942 191448 399122 191536
rect 399230 191448 399410 191536
rect 399518 191448 399698 191536
rect 399806 191448 399986 191536
rect 412286 191448 412466 191536
rect 412574 191448 412754 191536
rect 412862 191448 413042 191536
rect 413150 191448 413330 191536
rect 413438 191448 413618 191536
rect 413726 191448 413906 191536
rect 414014 191448 414194 191536
rect 414302 191448 414482 191536
rect 426782 191448 426962 191536
rect 427070 191448 427250 191536
rect 427358 191448 427538 191536
rect 427646 191448 427826 191536
rect 427934 191448 428114 191536
rect 428222 191448 428402 191536
rect 428510 191448 428690 191536
rect 428798 191448 428978 191536
rect 441278 191448 441458 191536
rect 441566 191448 441746 191536
rect 441854 191448 442034 191536
rect 442142 191448 442322 191536
rect 442430 191448 442610 191536
rect 442718 191448 442898 191536
rect 443006 191448 443186 191536
rect 443294 191448 443474 191536
rect 455774 191448 455954 191536
rect 456062 191448 456242 191536
rect 456350 191448 456530 191536
rect 456638 191448 456818 191536
rect 456926 191448 457106 191536
rect 457214 191448 457394 191536
rect 457502 191448 457682 191536
rect 457790 191448 457970 191536
rect 180350 191232 180530 191320
rect 180638 191232 180818 191320
rect 180926 191232 181106 191320
rect 181214 191232 181394 191320
rect 181502 191232 181682 191320
rect 181790 191232 181970 191320
rect 182078 191232 182258 191320
rect 182366 191232 182546 191320
rect 194846 191232 195026 191320
rect 195134 191232 195314 191320
rect 195422 191232 195602 191320
rect 195710 191232 195890 191320
rect 195998 191232 196178 191320
rect 196286 191232 196466 191320
rect 196574 191232 196754 191320
rect 196862 191232 197042 191320
rect 209342 191232 209522 191320
rect 209630 191232 209810 191320
rect 209918 191232 210098 191320
rect 210206 191232 210386 191320
rect 210494 191232 210674 191320
rect 210782 191232 210962 191320
rect 211070 191232 211250 191320
rect 211358 191232 211538 191320
rect 223838 191232 224018 191320
rect 224126 191232 224306 191320
rect 224414 191232 224594 191320
rect 224702 191232 224882 191320
rect 224990 191232 225170 191320
rect 225278 191232 225458 191320
rect 225566 191232 225746 191320
rect 225854 191232 226034 191320
rect 238334 191232 238514 191320
rect 238622 191232 238802 191320
rect 238910 191232 239090 191320
rect 239198 191232 239378 191320
rect 239486 191232 239666 191320
rect 239774 191232 239954 191320
rect 240062 191232 240242 191320
rect 240350 191232 240530 191320
rect 252830 191232 253010 191320
rect 253118 191232 253298 191320
rect 253406 191232 253586 191320
rect 253694 191232 253874 191320
rect 253982 191232 254162 191320
rect 254270 191232 254450 191320
rect 254558 191232 254738 191320
rect 254846 191232 255026 191320
rect 267326 191232 267506 191320
rect 267614 191232 267794 191320
rect 267902 191232 268082 191320
rect 268190 191232 268370 191320
rect 268478 191232 268658 191320
rect 268766 191232 268946 191320
rect 269054 191232 269234 191320
rect 269342 191232 269522 191320
rect 281822 191232 282002 191320
rect 282110 191232 282290 191320
rect 282398 191232 282578 191320
rect 282686 191232 282866 191320
rect 282974 191232 283154 191320
rect 283262 191232 283442 191320
rect 283550 191232 283730 191320
rect 283838 191232 284018 191320
rect 296318 191232 296498 191320
rect 296606 191232 296786 191320
rect 296894 191232 297074 191320
rect 297182 191232 297362 191320
rect 297470 191232 297650 191320
rect 297758 191232 297938 191320
rect 298046 191232 298226 191320
rect 298334 191232 298514 191320
rect 310814 191232 310994 191320
rect 311102 191232 311282 191320
rect 311390 191232 311570 191320
rect 311678 191232 311858 191320
rect 311966 191232 312146 191320
rect 312254 191232 312434 191320
rect 312542 191232 312722 191320
rect 312830 191232 313010 191320
rect 325310 191232 325490 191320
rect 325598 191232 325778 191320
rect 325886 191232 326066 191320
rect 326174 191232 326354 191320
rect 326462 191232 326642 191320
rect 326750 191232 326930 191320
rect 327038 191232 327218 191320
rect 327326 191232 327506 191320
rect 339806 191232 339986 191320
rect 340094 191232 340274 191320
rect 340382 191232 340562 191320
rect 340670 191232 340850 191320
rect 340958 191232 341138 191320
rect 341246 191232 341426 191320
rect 341534 191232 341714 191320
rect 341822 191232 342002 191320
rect 354302 191232 354482 191320
rect 354590 191232 354770 191320
rect 354878 191232 355058 191320
rect 355166 191232 355346 191320
rect 355454 191232 355634 191320
rect 355742 191232 355922 191320
rect 356030 191232 356210 191320
rect 356318 191232 356498 191320
rect 368798 191232 368978 191320
rect 369086 191232 369266 191320
rect 369374 191232 369554 191320
rect 369662 191232 369842 191320
rect 369950 191232 370130 191320
rect 370238 191232 370418 191320
rect 370526 191232 370706 191320
rect 370814 191232 370994 191320
rect 383294 191232 383474 191320
rect 383582 191232 383762 191320
rect 383870 191232 384050 191320
rect 384158 191232 384338 191320
rect 384446 191232 384626 191320
rect 384734 191232 384914 191320
rect 385022 191232 385202 191320
rect 385310 191232 385490 191320
rect 397790 191232 397970 191320
rect 398078 191232 398258 191320
rect 398366 191232 398546 191320
rect 398654 191232 398834 191320
rect 398942 191232 399122 191320
rect 399230 191232 399410 191320
rect 399518 191232 399698 191320
rect 399806 191232 399986 191320
rect 412286 191232 412466 191320
rect 412574 191232 412754 191320
rect 412862 191232 413042 191320
rect 413150 191232 413330 191320
rect 413438 191232 413618 191320
rect 413726 191232 413906 191320
rect 414014 191232 414194 191320
rect 414302 191232 414482 191320
rect 426782 191232 426962 191320
rect 427070 191232 427250 191320
rect 427358 191232 427538 191320
rect 427646 191232 427826 191320
rect 427934 191232 428114 191320
rect 428222 191232 428402 191320
rect 428510 191232 428690 191320
rect 428798 191232 428978 191320
rect 441278 191232 441458 191320
rect 441566 191232 441746 191320
rect 441854 191232 442034 191320
rect 442142 191232 442322 191320
rect 442430 191232 442610 191320
rect 442718 191232 442898 191320
rect 443006 191232 443186 191320
rect 443294 191232 443474 191320
rect 455774 191232 455954 191320
rect 456062 191232 456242 191320
rect 456350 191232 456530 191320
rect 456638 191232 456818 191320
rect 456926 191232 457106 191320
rect 457214 191232 457394 191320
rect 457502 191232 457682 191320
rect 457790 191232 457970 191320
rect 180350 190756 180530 190844
rect 180638 190756 180818 190844
rect 180926 190756 181106 190844
rect 181214 190756 181394 190844
rect 181502 190756 181682 190844
rect 181790 190756 181970 190844
rect 182078 190756 182258 190844
rect 182366 190756 182546 190844
rect 194846 190756 195026 190844
rect 195134 190756 195314 190844
rect 195422 190756 195602 190844
rect 195710 190756 195890 190844
rect 195998 190756 196178 190844
rect 196286 190756 196466 190844
rect 196574 190756 196754 190844
rect 196862 190756 197042 190844
rect 209342 190756 209522 190844
rect 209630 190756 209810 190844
rect 209918 190756 210098 190844
rect 210206 190756 210386 190844
rect 210494 190756 210674 190844
rect 210782 190756 210962 190844
rect 211070 190756 211250 190844
rect 211358 190756 211538 190844
rect 223838 190756 224018 190844
rect 224126 190756 224306 190844
rect 224414 190756 224594 190844
rect 224702 190756 224882 190844
rect 224990 190756 225170 190844
rect 225278 190756 225458 190844
rect 225566 190756 225746 190844
rect 225854 190756 226034 190844
rect 238334 190756 238514 190844
rect 238622 190756 238802 190844
rect 238910 190756 239090 190844
rect 239198 190756 239378 190844
rect 239486 190756 239666 190844
rect 239774 190756 239954 190844
rect 240062 190756 240242 190844
rect 240350 190756 240530 190844
rect 252830 190756 253010 190844
rect 253118 190756 253298 190844
rect 253406 190756 253586 190844
rect 253694 190756 253874 190844
rect 253982 190756 254162 190844
rect 254270 190756 254450 190844
rect 254558 190756 254738 190844
rect 254846 190756 255026 190844
rect 267326 190756 267506 190844
rect 267614 190756 267794 190844
rect 267902 190756 268082 190844
rect 268190 190756 268370 190844
rect 268478 190756 268658 190844
rect 268766 190756 268946 190844
rect 269054 190756 269234 190844
rect 269342 190756 269522 190844
rect 281822 190756 282002 190844
rect 282110 190756 282290 190844
rect 282398 190756 282578 190844
rect 282686 190756 282866 190844
rect 282974 190756 283154 190844
rect 283262 190756 283442 190844
rect 283550 190756 283730 190844
rect 283838 190756 284018 190844
rect 296318 190756 296498 190844
rect 296606 190756 296786 190844
rect 296894 190756 297074 190844
rect 297182 190756 297362 190844
rect 297470 190756 297650 190844
rect 297758 190756 297938 190844
rect 298046 190756 298226 190844
rect 298334 190756 298514 190844
rect 310814 190756 310994 190844
rect 311102 190756 311282 190844
rect 311390 190756 311570 190844
rect 311678 190756 311858 190844
rect 311966 190756 312146 190844
rect 312254 190756 312434 190844
rect 312542 190756 312722 190844
rect 312830 190756 313010 190844
rect 325310 190756 325490 190844
rect 325598 190756 325778 190844
rect 325886 190756 326066 190844
rect 326174 190756 326354 190844
rect 326462 190756 326642 190844
rect 326750 190756 326930 190844
rect 327038 190756 327218 190844
rect 327326 190756 327506 190844
rect 339806 190756 339986 190844
rect 340094 190756 340274 190844
rect 340382 190756 340562 190844
rect 340670 190756 340850 190844
rect 340958 190756 341138 190844
rect 341246 190756 341426 190844
rect 341534 190756 341714 190844
rect 341822 190756 342002 190844
rect 354302 190756 354482 190844
rect 354590 190756 354770 190844
rect 354878 190756 355058 190844
rect 355166 190756 355346 190844
rect 355454 190756 355634 190844
rect 355742 190756 355922 190844
rect 356030 190756 356210 190844
rect 356318 190756 356498 190844
rect 368798 190756 368978 190844
rect 369086 190756 369266 190844
rect 369374 190756 369554 190844
rect 369662 190756 369842 190844
rect 369950 190756 370130 190844
rect 370238 190756 370418 190844
rect 370526 190756 370706 190844
rect 370814 190756 370994 190844
rect 383294 190756 383474 190844
rect 383582 190756 383762 190844
rect 383870 190756 384050 190844
rect 384158 190756 384338 190844
rect 384446 190756 384626 190844
rect 384734 190756 384914 190844
rect 385022 190756 385202 190844
rect 385310 190756 385490 190844
rect 397790 190756 397970 190844
rect 398078 190756 398258 190844
rect 398366 190756 398546 190844
rect 398654 190756 398834 190844
rect 398942 190756 399122 190844
rect 399230 190756 399410 190844
rect 399518 190756 399698 190844
rect 399806 190756 399986 190844
rect 412286 190756 412466 190844
rect 412574 190756 412754 190844
rect 412862 190756 413042 190844
rect 413150 190756 413330 190844
rect 413438 190756 413618 190844
rect 413726 190756 413906 190844
rect 414014 190756 414194 190844
rect 414302 190756 414482 190844
rect 426782 190756 426962 190844
rect 427070 190756 427250 190844
rect 427358 190756 427538 190844
rect 427646 190756 427826 190844
rect 427934 190756 428114 190844
rect 428222 190756 428402 190844
rect 428510 190756 428690 190844
rect 428798 190756 428978 190844
rect 441278 190756 441458 190844
rect 441566 190756 441746 190844
rect 441854 190756 442034 190844
rect 442142 190756 442322 190844
rect 442430 190756 442610 190844
rect 442718 190756 442898 190844
rect 443006 190756 443186 190844
rect 443294 190756 443474 190844
rect 455774 190756 455954 190844
rect 456062 190756 456242 190844
rect 456350 190756 456530 190844
rect 456638 190756 456818 190844
rect 456926 190756 457106 190844
rect 457214 190756 457394 190844
rect 457502 190756 457682 190844
rect 457790 190756 457970 190844
rect 180350 190540 180530 190628
rect 180638 190540 180818 190628
rect 180926 190540 181106 190628
rect 181214 190540 181394 190628
rect 181502 190540 181682 190628
rect 181790 190540 181970 190628
rect 182078 190540 182258 190628
rect 182366 190540 182546 190628
rect 194846 190540 195026 190628
rect 195134 190540 195314 190628
rect 195422 190540 195602 190628
rect 195710 190540 195890 190628
rect 195998 190540 196178 190628
rect 196286 190540 196466 190628
rect 196574 190540 196754 190628
rect 196862 190540 197042 190628
rect 209342 190540 209522 190628
rect 209630 190540 209810 190628
rect 209918 190540 210098 190628
rect 210206 190540 210386 190628
rect 210494 190540 210674 190628
rect 210782 190540 210962 190628
rect 211070 190540 211250 190628
rect 211358 190540 211538 190628
rect 223838 190540 224018 190628
rect 224126 190540 224306 190628
rect 224414 190540 224594 190628
rect 224702 190540 224882 190628
rect 224990 190540 225170 190628
rect 225278 190540 225458 190628
rect 225566 190540 225746 190628
rect 225854 190540 226034 190628
rect 238334 190540 238514 190628
rect 238622 190540 238802 190628
rect 238910 190540 239090 190628
rect 239198 190540 239378 190628
rect 239486 190540 239666 190628
rect 239774 190540 239954 190628
rect 240062 190540 240242 190628
rect 240350 190540 240530 190628
rect 252830 190540 253010 190628
rect 253118 190540 253298 190628
rect 253406 190540 253586 190628
rect 253694 190540 253874 190628
rect 253982 190540 254162 190628
rect 254270 190540 254450 190628
rect 254558 190540 254738 190628
rect 254846 190540 255026 190628
rect 267326 190540 267506 190628
rect 267614 190540 267794 190628
rect 267902 190540 268082 190628
rect 268190 190540 268370 190628
rect 268478 190540 268658 190628
rect 268766 190540 268946 190628
rect 269054 190540 269234 190628
rect 269342 190540 269522 190628
rect 281822 190540 282002 190628
rect 282110 190540 282290 190628
rect 282398 190540 282578 190628
rect 282686 190540 282866 190628
rect 282974 190540 283154 190628
rect 283262 190540 283442 190628
rect 283550 190540 283730 190628
rect 283838 190540 284018 190628
rect 296318 190540 296498 190628
rect 296606 190540 296786 190628
rect 296894 190540 297074 190628
rect 297182 190540 297362 190628
rect 297470 190540 297650 190628
rect 297758 190540 297938 190628
rect 298046 190540 298226 190628
rect 298334 190540 298514 190628
rect 310814 190540 310994 190628
rect 311102 190540 311282 190628
rect 311390 190540 311570 190628
rect 311678 190540 311858 190628
rect 311966 190540 312146 190628
rect 312254 190540 312434 190628
rect 312542 190540 312722 190628
rect 312830 190540 313010 190628
rect 325310 190540 325490 190628
rect 325598 190540 325778 190628
rect 325886 190540 326066 190628
rect 326174 190540 326354 190628
rect 326462 190540 326642 190628
rect 326750 190540 326930 190628
rect 327038 190540 327218 190628
rect 327326 190540 327506 190628
rect 339806 190540 339986 190628
rect 340094 190540 340274 190628
rect 340382 190540 340562 190628
rect 340670 190540 340850 190628
rect 340958 190540 341138 190628
rect 341246 190540 341426 190628
rect 341534 190540 341714 190628
rect 341822 190540 342002 190628
rect 354302 190540 354482 190628
rect 354590 190540 354770 190628
rect 354878 190540 355058 190628
rect 355166 190540 355346 190628
rect 355454 190540 355634 190628
rect 355742 190540 355922 190628
rect 356030 190540 356210 190628
rect 356318 190540 356498 190628
rect 368798 190540 368978 190628
rect 369086 190540 369266 190628
rect 369374 190540 369554 190628
rect 369662 190540 369842 190628
rect 369950 190540 370130 190628
rect 370238 190540 370418 190628
rect 370526 190540 370706 190628
rect 370814 190540 370994 190628
rect 383294 190540 383474 190628
rect 383582 190540 383762 190628
rect 383870 190540 384050 190628
rect 384158 190540 384338 190628
rect 384446 190540 384626 190628
rect 384734 190540 384914 190628
rect 385022 190540 385202 190628
rect 385310 190540 385490 190628
rect 397790 190540 397970 190628
rect 398078 190540 398258 190628
rect 398366 190540 398546 190628
rect 398654 190540 398834 190628
rect 398942 190540 399122 190628
rect 399230 190540 399410 190628
rect 399518 190540 399698 190628
rect 399806 190540 399986 190628
rect 412286 190540 412466 190628
rect 412574 190540 412754 190628
rect 412862 190540 413042 190628
rect 413150 190540 413330 190628
rect 413438 190540 413618 190628
rect 413726 190540 413906 190628
rect 414014 190540 414194 190628
rect 414302 190540 414482 190628
rect 426782 190540 426962 190628
rect 427070 190540 427250 190628
rect 427358 190540 427538 190628
rect 427646 190540 427826 190628
rect 427934 190540 428114 190628
rect 428222 190540 428402 190628
rect 428510 190540 428690 190628
rect 428798 190540 428978 190628
rect 441278 190540 441458 190628
rect 441566 190540 441746 190628
rect 441854 190540 442034 190628
rect 442142 190540 442322 190628
rect 442430 190540 442610 190628
rect 442718 190540 442898 190628
rect 443006 190540 443186 190628
rect 443294 190540 443474 190628
rect 455774 190540 455954 190628
rect 456062 190540 456242 190628
rect 456350 190540 456530 190628
rect 456638 190540 456818 190628
rect 456926 190540 457106 190628
rect 457214 190540 457394 190628
rect 457502 190540 457682 190628
rect 457790 190540 457970 190628
rect 180350 176388 180530 176476
rect 180638 176388 180818 176476
rect 180926 176388 181106 176476
rect 181214 176388 181394 176476
rect 181502 176388 181682 176476
rect 181790 176388 181970 176476
rect 182078 176388 182258 176476
rect 182366 176388 182546 176476
rect 194846 176388 195026 176476
rect 195134 176388 195314 176476
rect 195422 176388 195602 176476
rect 195710 176388 195890 176476
rect 195998 176388 196178 176476
rect 196286 176388 196466 176476
rect 196574 176388 196754 176476
rect 196862 176388 197042 176476
rect 209342 176388 209522 176476
rect 209630 176388 209810 176476
rect 209918 176388 210098 176476
rect 210206 176388 210386 176476
rect 210494 176388 210674 176476
rect 210782 176388 210962 176476
rect 211070 176388 211250 176476
rect 211358 176388 211538 176476
rect 223838 176388 224018 176476
rect 224126 176388 224306 176476
rect 224414 176388 224594 176476
rect 224702 176388 224882 176476
rect 224990 176388 225170 176476
rect 225278 176388 225458 176476
rect 225566 176388 225746 176476
rect 225854 176388 226034 176476
rect 238334 176388 238514 176476
rect 238622 176388 238802 176476
rect 238910 176388 239090 176476
rect 239198 176388 239378 176476
rect 239486 176388 239666 176476
rect 239774 176388 239954 176476
rect 240062 176388 240242 176476
rect 240350 176388 240530 176476
rect 252830 176388 253010 176476
rect 253118 176388 253298 176476
rect 253406 176388 253586 176476
rect 253694 176388 253874 176476
rect 253982 176388 254162 176476
rect 254270 176388 254450 176476
rect 254558 176388 254738 176476
rect 254846 176388 255026 176476
rect 267326 176388 267506 176476
rect 267614 176388 267794 176476
rect 267902 176388 268082 176476
rect 268190 176388 268370 176476
rect 268478 176388 268658 176476
rect 268766 176388 268946 176476
rect 269054 176388 269234 176476
rect 269342 176388 269522 176476
rect 281822 176388 282002 176476
rect 282110 176388 282290 176476
rect 282398 176388 282578 176476
rect 282686 176388 282866 176476
rect 282974 176388 283154 176476
rect 283262 176388 283442 176476
rect 283550 176388 283730 176476
rect 283838 176388 284018 176476
rect 296318 176388 296498 176476
rect 296606 176388 296786 176476
rect 296894 176388 297074 176476
rect 297182 176388 297362 176476
rect 297470 176388 297650 176476
rect 297758 176388 297938 176476
rect 298046 176388 298226 176476
rect 298334 176388 298514 176476
rect 310814 176388 310994 176476
rect 311102 176388 311282 176476
rect 311390 176388 311570 176476
rect 311678 176388 311858 176476
rect 311966 176388 312146 176476
rect 312254 176388 312434 176476
rect 312542 176388 312722 176476
rect 312830 176388 313010 176476
rect 325310 176388 325490 176476
rect 325598 176388 325778 176476
rect 325886 176388 326066 176476
rect 326174 176388 326354 176476
rect 326462 176388 326642 176476
rect 326750 176388 326930 176476
rect 327038 176388 327218 176476
rect 327326 176388 327506 176476
rect 339806 176388 339986 176476
rect 340094 176388 340274 176476
rect 340382 176388 340562 176476
rect 340670 176388 340850 176476
rect 340958 176388 341138 176476
rect 341246 176388 341426 176476
rect 341534 176388 341714 176476
rect 341822 176388 342002 176476
rect 354302 176388 354482 176476
rect 354590 176388 354770 176476
rect 354878 176388 355058 176476
rect 355166 176388 355346 176476
rect 355454 176388 355634 176476
rect 355742 176388 355922 176476
rect 356030 176388 356210 176476
rect 356318 176388 356498 176476
rect 368798 176388 368978 176476
rect 369086 176388 369266 176476
rect 369374 176388 369554 176476
rect 369662 176388 369842 176476
rect 369950 176388 370130 176476
rect 370238 176388 370418 176476
rect 370526 176388 370706 176476
rect 370814 176388 370994 176476
rect 383294 176388 383474 176476
rect 383582 176388 383762 176476
rect 383870 176388 384050 176476
rect 384158 176388 384338 176476
rect 384446 176388 384626 176476
rect 384734 176388 384914 176476
rect 385022 176388 385202 176476
rect 385310 176388 385490 176476
rect 397790 176388 397970 176476
rect 398078 176388 398258 176476
rect 398366 176388 398546 176476
rect 398654 176388 398834 176476
rect 398942 176388 399122 176476
rect 399230 176388 399410 176476
rect 399518 176388 399698 176476
rect 399806 176388 399986 176476
rect 412286 176388 412466 176476
rect 412574 176388 412754 176476
rect 412862 176388 413042 176476
rect 413150 176388 413330 176476
rect 413438 176388 413618 176476
rect 413726 176388 413906 176476
rect 414014 176388 414194 176476
rect 414302 176388 414482 176476
rect 426782 176388 426962 176476
rect 427070 176388 427250 176476
rect 427358 176388 427538 176476
rect 427646 176388 427826 176476
rect 427934 176388 428114 176476
rect 428222 176388 428402 176476
rect 428510 176388 428690 176476
rect 428798 176388 428978 176476
rect 441278 176388 441458 176476
rect 441566 176388 441746 176476
rect 441854 176388 442034 176476
rect 442142 176388 442322 176476
rect 442430 176388 442610 176476
rect 442718 176388 442898 176476
rect 443006 176388 443186 176476
rect 443294 176388 443474 176476
rect 455774 176388 455954 176476
rect 456062 176388 456242 176476
rect 456350 176388 456530 176476
rect 456638 176388 456818 176476
rect 456926 176388 457106 176476
rect 457214 176388 457394 176476
rect 457502 176388 457682 176476
rect 457790 176388 457970 176476
rect 180350 176172 180530 176260
rect 180638 176172 180818 176260
rect 180926 176172 181106 176260
rect 181214 176172 181394 176260
rect 181502 176172 181682 176260
rect 181790 176172 181970 176260
rect 182078 176172 182258 176260
rect 182366 176172 182546 176260
rect 194846 176172 195026 176260
rect 195134 176172 195314 176260
rect 195422 176172 195602 176260
rect 195710 176172 195890 176260
rect 195998 176172 196178 176260
rect 196286 176172 196466 176260
rect 196574 176172 196754 176260
rect 196862 176172 197042 176260
rect 209342 176172 209522 176260
rect 209630 176172 209810 176260
rect 209918 176172 210098 176260
rect 210206 176172 210386 176260
rect 210494 176172 210674 176260
rect 210782 176172 210962 176260
rect 211070 176172 211250 176260
rect 211358 176172 211538 176260
rect 223838 176172 224018 176260
rect 224126 176172 224306 176260
rect 224414 176172 224594 176260
rect 224702 176172 224882 176260
rect 224990 176172 225170 176260
rect 225278 176172 225458 176260
rect 225566 176172 225746 176260
rect 225854 176172 226034 176260
rect 238334 176172 238514 176260
rect 238622 176172 238802 176260
rect 238910 176172 239090 176260
rect 239198 176172 239378 176260
rect 239486 176172 239666 176260
rect 239774 176172 239954 176260
rect 240062 176172 240242 176260
rect 240350 176172 240530 176260
rect 252830 176172 253010 176260
rect 253118 176172 253298 176260
rect 253406 176172 253586 176260
rect 253694 176172 253874 176260
rect 253982 176172 254162 176260
rect 254270 176172 254450 176260
rect 254558 176172 254738 176260
rect 254846 176172 255026 176260
rect 267326 176172 267506 176260
rect 267614 176172 267794 176260
rect 267902 176172 268082 176260
rect 268190 176172 268370 176260
rect 268478 176172 268658 176260
rect 268766 176172 268946 176260
rect 269054 176172 269234 176260
rect 269342 176172 269522 176260
rect 281822 176172 282002 176260
rect 282110 176172 282290 176260
rect 282398 176172 282578 176260
rect 282686 176172 282866 176260
rect 282974 176172 283154 176260
rect 283262 176172 283442 176260
rect 283550 176172 283730 176260
rect 283838 176172 284018 176260
rect 296318 176172 296498 176260
rect 296606 176172 296786 176260
rect 296894 176172 297074 176260
rect 297182 176172 297362 176260
rect 297470 176172 297650 176260
rect 297758 176172 297938 176260
rect 298046 176172 298226 176260
rect 298334 176172 298514 176260
rect 310814 176172 310994 176260
rect 311102 176172 311282 176260
rect 311390 176172 311570 176260
rect 311678 176172 311858 176260
rect 311966 176172 312146 176260
rect 312254 176172 312434 176260
rect 312542 176172 312722 176260
rect 312830 176172 313010 176260
rect 325310 176172 325490 176260
rect 325598 176172 325778 176260
rect 325886 176172 326066 176260
rect 326174 176172 326354 176260
rect 326462 176172 326642 176260
rect 326750 176172 326930 176260
rect 327038 176172 327218 176260
rect 327326 176172 327506 176260
rect 339806 176172 339986 176260
rect 340094 176172 340274 176260
rect 340382 176172 340562 176260
rect 340670 176172 340850 176260
rect 340958 176172 341138 176260
rect 341246 176172 341426 176260
rect 341534 176172 341714 176260
rect 341822 176172 342002 176260
rect 354302 176172 354482 176260
rect 354590 176172 354770 176260
rect 354878 176172 355058 176260
rect 355166 176172 355346 176260
rect 355454 176172 355634 176260
rect 355742 176172 355922 176260
rect 356030 176172 356210 176260
rect 356318 176172 356498 176260
rect 368798 176172 368978 176260
rect 369086 176172 369266 176260
rect 369374 176172 369554 176260
rect 369662 176172 369842 176260
rect 369950 176172 370130 176260
rect 370238 176172 370418 176260
rect 370526 176172 370706 176260
rect 370814 176172 370994 176260
rect 383294 176172 383474 176260
rect 383582 176172 383762 176260
rect 383870 176172 384050 176260
rect 384158 176172 384338 176260
rect 384446 176172 384626 176260
rect 384734 176172 384914 176260
rect 385022 176172 385202 176260
rect 385310 176172 385490 176260
rect 397790 176172 397970 176260
rect 398078 176172 398258 176260
rect 398366 176172 398546 176260
rect 398654 176172 398834 176260
rect 398942 176172 399122 176260
rect 399230 176172 399410 176260
rect 399518 176172 399698 176260
rect 399806 176172 399986 176260
rect 412286 176172 412466 176260
rect 412574 176172 412754 176260
rect 412862 176172 413042 176260
rect 413150 176172 413330 176260
rect 413438 176172 413618 176260
rect 413726 176172 413906 176260
rect 414014 176172 414194 176260
rect 414302 176172 414482 176260
rect 426782 176172 426962 176260
rect 427070 176172 427250 176260
rect 427358 176172 427538 176260
rect 427646 176172 427826 176260
rect 427934 176172 428114 176260
rect 428222 176172 428402 176260
rect 428510 176172 428690 176260
rect 428798 176172 428978 176260
rect 441278 176172 441458 176260
rect 441566 176172 441746 176260
rect 441854 176172 442034 176260
rect 442142 176172 442322 176260
rect 442430 176172 442610 176260
rect 442718 176172 442898 176260
rect 443006 176172 443186 176260
rect 443294 176172 443474 176260
rect 455774 176172 455954 176260
rect 456062 176172 456242 176260
rect 456350 176172 456530 176260
rect 456638 176172 456818 176260
rect 456926 176172 457106 176260
rect 457214 176172 457394 176260
rect 457502 176172 457682 176260
rect 457790 176172 457970 176260
rect 180350 175696 180530 175784
rect 180638 175696 180818 175784
rect 180926 175696 181106 175784
rect 181214 175696 181394 175784
rect 181502 175696 181682 175784
rect 181790 175696 181970 175784
rect 182078 175696 182258 175784
rect 182366 175696 182546 175784
rect 194846 175696 195026 175784
rect 195134 175696 195314 175784
rect 195422 175696 195602 175784
rect 195710 175696 195890 175784
rect 195998 175696 196178 175784
rect 196286 175696 196466 175784
rect 196574 175696 196754 175784
rect 196862 175696 197042 175784
rect 209342 175696 209522 175784
rect 209630 175696 209810 175784
rect 209918 175696 210098 175784
rect 210206 175696 210386 175784
rect 210494 175696 210674 175784
rect 210782 175696 210962 175784
rect 211070 175696 211250 175784
rect 211358 175696 211538 175784
rect 223838 175696 224018 175784
rect 224126 175696 224306 175784
rect 224414 175696 224594 175784
rect 224702 175696 224882 175784
rect 224990 175696 225170 175784
rect 225278 175696 225458 175784
rect 225566 175696 225746 175784
rect 225854 175696 226034 175784
rect 238334 175696 238514 175784
rect 238622 175696 238802 175784
rect 238910 175696 239090 175784
rect 239198 175696 239378 175784
rect 239486 175696 239666 175784
rect 239774 175696 239954 175784
rect 240062 175696 240242 175784
rect 240350 175696 240530 175784
rect 252830 175696 253010 175784
rect 253118 175696 253298 175784
rect 253406 175696 253586 175784
rect 253694 175696 253874 175784
rect 253982 175696 254162 175784
rect 254270 175696 254450 175784
rect 254558 175696 254738 175784
rect 254846 175696 255026 175784
rect 267326 175696 267506 175784
rect 267614 175696 267794 175784
rect 267902 175696 268082 175784
rect 268190 175696 268370 175784
rect 268478 175696 268658 175784
rect 268766 175696 268946 175784
rect 269054 175696 269234 175784
rect 269342 175696 269522 175784
rect 281822 175696 282002 175784
rect 282110 175696 282290 175784
rect 282398 175696 282578 175784
rect 282686 175696 282866 175784
rect 282974 175696 283154 175784
rect 283262 175696 283442 175784
rect 283550 175696 283730 175784
rect 283838 175696 284018 175784
rect 296318 175696 296498 175784
rect 296606 175696 296786 175784
rect 296894 175696 297074 175784
rect 297182 175696 297362 175784
rect 297470 175696 297650 175784
rect 297758 175696 297938 175784
rect 298046 175696 298226 175784
rect 298334 175696 298514 175784
rect 310814 175696 310994 175784
rect 311102 175696 311282 175784
rect 311390 175696 311570 175784
rect 311678 175696 311858 175784
rect 311966 175696 312146 175784
rect 312254 175696 312434 175784
rect 312542 175696 312722 175784
rect 312830 175696 313010 175784
rect 325310 175696 325490 175784
rect 325598 175696 325778 175784
rect 325886 175696 326066 175784
rect 326174 175696 326354 175784
rect 326462 175696 326642 175784
rect 326750 175696 326930 175784
rect 327038 175696 327218 175784
rect 327326 175696 327506 175784
rect 339806 175696 339986 175784
rect 340094 175696 340274 175784
rect 340382 175696 340562 175784
rect 340670 175696 340850 175784
rect 340958 175696 341138 175784
rect 341246 175696 341426 175784
rect 341534 175696 341714 175784
rect 341822 175696 342002 175784
rect 354302 175696 354482 175784
rect 354590 175696 354770 175784
rect 354878 175696 355058 175784
rect 355166 175696 355346 175784
rect 355454 175696 355634 175784
rect 355742 175696 355922 175784
rect 356030 175696 356210 175784
rect 356318 175696 356498 175784
rect 368798 175696 368978 175784
rect 369086 175696 369266 175784
rect 369374 175696 369554 175784
rect 369662 175696 369842 175784
rect 369950 175696 370130 175784
rect 370238 175696 370418 175784
rect 370526 175696 370706 175784
rect 370814 175696 370994 175784
rect 383294 175696 383474 175784
rect 383582 175696 383762 175784
rect 383870 175696 384050 175784
rect 384158 175696 384338 175784
rect 384446 175696 384626 175784
rect 384734 175696 384914 175784
rect 385022 175696 385202 175784
rect 385310 175696 385490 175784
rect 397790 175696 397970 175784
rect 398078 175696 398258 175784
rect 398366 175696 398546 175784
rect 398654 175696 398834 175784
rect 398942 175696 399122 175784
rect 399230 175696 399410 175784
rect 399518 175696 399698 175784
rect 399806 175696 399986 175784
rect 412286 175696 412466 175784
rect 412574 175696 412754 175784
rect 412862 175696 413042 175784
rect 413150 175696 413330 175784
rect 413438 175696 413618 175784
rect 413726 175696 413906 175784
rect 414014 175696 414194 175784
rect 414302 175696 414482 175784
rect 426782 175696 426962 175784
rect 427070 175696 427250 175784
rect 427358 175696 427538 175784
rect 427646 175696 427826 175784
rect 427934 175696 428114 175784
rect 428222 175696 428402 175784
rect 428510 175696 428690 175784
rect 428798 175696 428978 175784
rect 441278 175696 441458 175784
rect 441566 175696 441746 175784
rect 441854 175696 442034 175784
rect 442142 175696 442322 175784
rect 442430 175696 442610 175784
rect 442718 175696 442898 175784
rect 443006 175696 443186 175784
rect 443294 175696 443474 175784
rect 455774 175696 455954 175784
rect 456062 175696 456242 175784
rect 456350 175696 456530 175784
rect 456638 175696 456818 175784
rect 456926 175696 457106 175784
rect 457214 175696 457394 175784
rect 457502 175696 457682 175784
rect 457790 175696 457970 175784
rect 180350 175480 180530 175568
rect 180638 175480 180818 175568
rect 180926 175480 181106 175568
rect 181214 175480 181394 175568
rect 181502 175480 181682 175568
rect 181790 175480 181970 175568
rect 182078 175480 182258 175568
rect 182366 175480 182546 175568
rect 194846 175480 195026 175568
rect 195134 175480 195314 175568
rect 195422 175480 195602 175568
rect 195710 175480 195890 175568
rect 195998 175480 196178 175568
rect 196286 175480 196466 175568
rect 196574 175480 196754 175568
rect 196862 175480 197042 175568
rect 209342 175480 209522 175568
rect 209630 175480 209810 175568
rect 209918 175480 210098 175568
rect 210206 175480 210386 175568
rect 210494 175480 210674 175568
rect 210782 175480 210962 175568
rect 211070 175480 211250 175568
rect 211358 175480 211538 175568
rect 223838 175480 224018 175568
rect 224126 175480 224306 175568
rect 224414 175480 224594 175568
rect 224702 175480 224882 175568
rect 224990 175480 225170 175568
rect 225278 175480 225458 175568
rect 225566 175480 225746 175568
rect 225854 175480 226034 175568
rect 238334 175480 238514 175568
rect 238622 175480 238802 175568
rect 238910 175480 239090 175568
rect 239198 175480 239378 175568
rect 239486 175480 239666 175568
rect 239774 175480 239954 175568
rect 240062 175480 240242 175568
rect 240350 175480 240530 175568
rect 252830 175480 253010 175568
rect 253118 175480 253298 175568
rect 253406 175480 253586 175568
rect 253694 175480 253874 175568
rect 253982 175480 254162 175568
rect 254270 175480 254450 175568
rect 254558 175480 254738 175568
rect 254846 175480 255026 175568
rect 267326 175480 267506 175568
rect 267614 175480 267794 175568
rect 267902 175480 268082 175568
rect 268190 175480 268370 175568
rect 268478 175480 268658 175568
rect 268766 175480 268946 175568
rect 269054 175480 269234 175568
rect 269342 175480 269522 175568
rect 281822 175480 282002 175568
rect 282110 175480 282290 175568
rect 282398 175480 282578 175568
rect 282686 175480 282866 175568
rect 282974 175480 283154 175568
rect 283262 175480 283442 175568
rect 283550 175480 283730 175568
rect 283838 175480 284018 175568
rect 296318 175480 296498 175568
rect 296606 175480 296786 175568
rect 296894 175480 297074 175568
rect 297182 175480 297362 175568
rect 297470 175480 297650 175568
rect 297758 175480 297938 175568
rect 298046 175480 298226 175568
rect 298334 175480 298514 175568
rect 310814 175480 310994 175568
rect 311102 175480 311282 175568
rect 311390 175480 311570 175568
rect 311678 175480 311858 175568
rect 311966 175480 312146 175568
rect 312254 175480 312434 175568
rect 312542 175480 312722 175568
rect 312830 175480 313010 175568
rect 325310 175480 325490 175568
rect 325598 175480 325778 175568
rect 325886 175480 326066 175568
rect 326174 175480 326354 175568
rect 326462 175480 326642 175568
rect 326750 175480 326930 175568
rect 327038 175480 327218 175568
rect 327326 175480 327506 175568
rect 339806 175480 339986 175568
rect 340094 175480 340274 175568
rect 340382 175480 340562 175568
rect 340670 175480 340850 175568
rect 340958 175480 341138 175568
rect 341246 175480 341426 175568
rect 341534 175480 341714 175568
rect 341822 175480 342002 175568
rect 354302 175480 354482 175568
rect 354590 175480 354770 175568
rect 354878 175480 355058 175568
rect 355166 175480 355346 175568
rect 355454 175480 355634 175568
rect 355742 175480 355922 175568
rect 356030 175480 356210 175568
rect 356318 175480 356498 175568
rect 368798 175480 368978 175568
rect 369086 175480 369266 175568
rect 369374 175480 369554 175568
rect 369662 175480 369842 175568
rect 369950 175480 370130 175568
rect 370238 175480 370418 175568
rect 370526 175480 370706 175568
rect 370814 175480 370994 175568
rect 383294 175480 383474 175568
rect 383582 175480 383762 175568
rect 383870 175480 384050 175568
rect 384158 175480 384338 175568
rect 384446 175480 384626 175568
rect 384734 175480 384914 175568
rect 385022 175480 385202 175568
rect 385310 175480 385490 175568
rect 397790 175480 397970 175568
rect 398078 175480 398258 175568
rect 398366 175480 398546 175568
rect 398654 175480 398834 175568
rect 398942 175480 399122 175568
rect 399230 175480 399410 175568
rect 399518 175480 399698 175568
rect 399806 175480 399986 175568
rect 412286 175480 412466 175568
rect 412574 175480 412754 175568
rect 412862 175480 413042 175568
rect 413150 175480 413330 175568
rect 413438 175480 413618 175568
rect 413726 175480 413906 175568
rect 414014 175480 414194 175568
rect 414302 175480 414482 175568
rect 426782 175480 426962 175568
rect 427070 175480 427250 175568
rect 427358 175480 427538 175568
rect 427646 175480 427826 175568
rect 427934 175480 428114 175568
rect 428222 175480 428402 175568
rect 428510 175480 428690 175568
rect 428798 175480 428978 175568
rect 441278 175480 441458 175568
rect 441566 175480 441746 175568
rect 441854 175480 442034 175568
rect 442142 175480 442322 175568
rect 442430 175480 442610 175568
rect 442718 175480 442898 175568
rect 443006 175480 443186 175568
rect 443294 175480 443474 175568
rect 455774 175480 455954 175568
rect 456062 175480 456242 175568
rect 456350 175480 456530 175568
rect 456638 175480 456818 175568
rect 456926 175480 457106 175568
rect 457214 175480 457394 175568
rect 457502 175480 457682 175568
rect 457790 175480 457970 175568
rect 180350 161328 180530 161416
rect 180638 161328 180818 161416
rect 180926 161328 181106 161416
rect 181214 161328 181394 161416
rect 181502 161328 181682 161416
rect 181790 161328 181970 161416
rect 182078 161328 182258 161416
rect 182366 161328 182546 161416
rect 194846 161328 195026 161416
rect 195134 161328 195314 161416
rect 195422 161328 195602 161416
rect 195710 161328 195890 161416
rect 195998 161328 196178 161416
rect 196286 161328 196466 161416
rect 196574 161328 196754 161416
rect 196862 161328 197042 161416
rect 209342 161328 209522 161416
rect 209630 161328 209810 161416
rect 209918 161328 210098 161416
rect 210206 161328 210386 161416
rect 210494 161328 210674 161416
rect 210782 161328 210962 161416
rect 211070 161328 211250 161416
rect 211358 161328 211538 161416
rect 223838 161328 224018 161416
rect 224126 161328 224306 161416
rect 224414 161328 224594 161416
rect 224702 161328 224882 161416
rect 224990 161328 225170 161416
rect 225278 161328 225458 161416
rect 225566 161328 225746 161416
rect 225854 161328 226034 161416
rect 238334 161328 238514 161416
rect 238622 161328 238802 161416
rect 238910 161328 239090 161416
rect 239198 161328 239378 161416
rect 239486 161328 239666 161416
rect 239774 161328 239954 161416
rect 240062 161328 240242 161416
rect 240350 161328 240530 161416
rect 252830 161328 253010 161416
rect 253118 161328 253298 161416
rect 253406 161328 253586 161416
rect 253694 161328 253874 161416
rect 253982 161328 254162 161416
rect 254270 161328 254450 161416
rect 254558 161328 254738 161416
rect 254846 161328 255026 161416
rect 267326 161328 267506 161416
rect 267614 161328 267794 161416
rect 267902 161328 268082 161416
rect 268190 161328 268370 161416
rect 268478 161328 268658 161416
rect 268766 161328 268946 161416
rect 269054 161328 269234 161416
rect 269342 161328 269522 161416
rect 281822 161328 282002 161416
rect 282110 161328 282290 161416
rect 282398 161328 282578 161416
rect 282686 161328 282866 161416
rect 282974 161328 283154 161416
rect 283262 161328 283442 161416
rect 283550 161328 283730 161416
rect 283838 161328 284018 161416
rect 296318 161328 296498 161416
rect 296606 161328 296786 161416
rect 296894 161328 297074 161416
rect 297182 161328 297362 161416
rect 297470 161328 297650 161416
rect 297758 161328 297938 161416
rect 298046 161328 298226 161416
rect 298334 161328 298514 161416
rect 310814 161328 310994 161416
rect 311102 161328 311282 161416
rect 311390 161328 311570 161416
rect 311678 161328 311858 161416
rect 311966 161328 312146 161416
rect 312254 161328 312434 161416
rect 312542 161328 312722 161416
rect 312830 161328 313010 161416
rect 325310 161328 325490 161416
rect 325598 161328 325778 161416
rect 325886 161328 326066 161416
rect 326174 161328 326354 161416
rect 326462 161328 326642 161416
rect 326750 161328 326930 161416
rect 327038 161328 327218 161416
rect 327326 161328 327506 161416
rect 339806 161328 339986 161416
rect 340094 161328 340274 161416
rect 340382 161328 340562 161416
rect 340670 161328 340850 161416
rect 340958 161328 341138 161416
rect 341246 161328 341426 161416
rect 341534 161328 341714 161416
rect 341822 161328 342002 161416
rect 354302 161328 354482 161416
rect 354590 161328 354770 161416
rect 354878 161328 355058 161416
rect 355166 161328 355346 161416
rect 355454 161328 355634 161416
rect 355742 161328 355922 161416
rect 356030 161328 356210 161416
rect 356318 161328 356498 161416
rect 368798 161328 368978 161416
rect 369086 161328 369266 161416
rect 369374 161328 369554 161416
rect 369662 161328 369842 161416
rect 369950 161328 370130 161416
rect 370238 161328 370418 161416
rect 370526 161328 370706 161416
rect 370814 161328 370994 161416
rect 383294 161328 383474 161416
rect 383582 161328 383762 161416
rect 383870 161328 384050 161416
rect 384158 161328 384338 161416
rect 384446 161328 384626 161416
rect 384734 161328 384914 161416
rect 385022 161328 385202 161416
rect 385310 161328 385490 161416
rect 397790 161328 397970 161416
rect 398078 161328 398258 161416
rect 398366 161328 398546 161416
rect 398654 161328 398834 161416
rect 398942 161328 399122 161416
rect 399230 161328 399410 161416
rect 399518 161328 399698 161416
rect 399806 161328 399986 161416
rect 412286 161328 412466 161416
rect 412574 161328 412754 161416
rect 412862 161328 413042 161416
rect 413150 161328 413330 161416
rect 413438 161328 413618 161416
rect 413726 161328 413906 161416
rect 414014 161328 414194 161416
rect 414302 161328 414482 161416
rect 426782 161328 426962 161416
rect 427070 161328 427250 161416
rect 427358 161328 427538 161416
rect 427646 161328 427826 161416
rect 427934 161328 428114 161416
rect 428222 161328 428402 161416
rect 428510 161328 428690 161416
rect 428798 161328 428978 161416
rect 441278 161328 441458 161416
rect 441566 161328 441746 161416
rect 441854 161328 442034 161416
rect 442142 161328 442322 161416
rect 442430 161328 442610 161416
rect 442718 161328 442898 161416
rect 443006 161328 443186 161416
rect 443294 161328 443474 161416
rect 455774 161328 455954 161416
rect 456062 161328 456242 161416
rect 456350 161328 456530 161416
rect 456638 161328 456818 161416
rect 456926 161328 457106 161416
rect 457214 161328 457394 161416
rect 457502 161328 457682 161416
rect 457790 161328 457970 161416
rect 180350 161112 180530 161200
rect 180638 161112 180818 161200
rect 180926 161112 181106 161200
rect 181214 161112 181394 161200
rect 181502 161112 181682 161200
rect 181790 161112 181970 161200
rect 182078 161112 182258 161200
rect 182366 161112 182546 161200
rect 194846 161112 195026 161200
rect 195134 161112 195314 161200
rect 195422 161112 195602 161200
rect 195710 161112 195890 161200
rect 195998 161112 196178 161200
rect 196286 161112 196466 161200
rect 196574 161112 196754 161200
rect 196862 161112 197042 161200
rect 209342 161112 209522 161200
rect 209630 161112 209810 161200
rect 209918 161112 210098 161200
rect 210206 161112 210386 161200
rect 210494 161112 210674 161200
rect 210782 161112 210962 161200
rect 211070 161112 211250 161200
rect 211358 161112 211538 161200
rect 223838 161112 224018 161200
rect 224126 161112 224306 161200
rect 224414 161112 224594 161200
rect 224702 161112 224882 161200
rect 224990 161112 225170 161200
rect 225278 161112 225458 161200
rect 225566 161112 225746 161200
rect 225854 161112 226034 161200
rect 238334 161112 238514 161200
rect 238622 161112 238802 161200
rect 238910 161112 239090 161200
rect 239198 161112 239378 161200
rect 239486 161112 239666 161200
rect 239774 161112 239954 161200
rect 240062 161112 240242 161200
rect 240350 161112 240530 161200
rect 252830 161112 253010 161200
rect 253118 161112 253298 161200
rect 253406 161112 253586 161200
rect 253694 161112 253874 161200
rect 253982 161112 254162 161200
rect 254270 161112 254450 161200
rect 254558 161112 254738 161200
rect 254846 161112 255026 161200
rect 267326 161112 267506 161200
rect 267614 161112 267794 161200
rect 267902 161112 268082 161200
rect 268190 161112 268370 161200
rect 268478 161112 268658 161200
rect 268766 161112 268946 161200
rect 269054 161112 269234 161200
rect 269342 161112 269522 161200
rect 281822 161112 282002 161200
rect 282110 161112 282290 161200
rect 282398 161112 282578 161200
rect 282686 161112 282866 161200
rect 282974 161112 283154 161200
rect 283262 161112 283442 161200
rect 283550 161112 283730 161200
rect 283838 161112 284018 161200
rect 296318 161112 296498 161200
rect 296606 161112 296786 161200
rect 296894 161112 297074 161200
rect 297182 161112 297362 161200
rect 297470 161112 297650 161200
rect 297758 161112 297938 161200
rect 298046 161112 298226 161200
rect 298334 161112 298514 161200
rect 310814 161112 310994 161200
rect 311102 161112 311282 161200
rect 311390 161112 311570 161200
rect 311678 161112 311858 161200
rect 311966 161112 312146 161200
rect 312254 161112 312434 161200
rect 312542 161112 312722 161200
rect 312830 161112 313010 161200
rect 325310 161112 325490 161200
rect 325598 161112 325778 161200
rect 325886 161112 326066 161200
rect 326174 161112 326354 161200
rect 326462 161112 326642 161200
rect 326750 161112 326930 161200
rect 327038 161112 327218 161200
rect 327326 161112 327506 161200
rect 339806 161112 339986 161200
rect 340094 161112 340274 161200
rect 340382 161112 340562 161200
rect 340670 161112 340850 161200
rect 340958 161112 341138 161200
rect 341246 161112 341426 161200
rect 341534 161112 341714 161200
rect 341822 161112 342002 161200
rect 354302 161112 354482 161200
rect 354590 161112 354770 161200
rect 354878 161112 355058 161200
rect 355166 161112 355346 161200
rect 355454 161112 355634 161200
rect 355742 161112 355922 161200
rect 356030 161112 356210 161200
rect 356318 161112 356498 161200
rect 368798 161112 368978 161200
rect 369086 161112 369266 161200
rect 369374 161112 369554 161200
rect 369662 161112 369842 161200
rect 369950 161112 370130 161200
rect 370238 161112 370418 161200
rect 370526 161112 370706 161200
rect 370814 161112 370994 161200
rect 383294 161112 383474 161200
rect 383582 161112 383762 161200
rect 383870 161112 384050 161200
rect 384158 161112 384338 161200
rect 384446 161112 384626 161200
rect 384734 161112 384914 161200
rect 385022 161112 385202 161200
rect 385310 161112 385490 161200
rect 397790 161112 397970 161200
rect 398078 161112 398258 161200
rect 398366 161112 398546 161200
rect 398654 161112 398834 161200
rect 398942 161112 399122 161200
rect 399230 161112 399410 161200
rect 399518 161112 399698 161200
rect 399806 161112 399986 161200
rect 412286 161112 412466 161200
rect 412574 161112 412754 161200
rect 412862 161112 413042 161200
rect 413150 161112 413330 161200
rect 413438 161112 413618 161200
rect 413726 161112 413906 161200
rect 414014 161112 414194 161200
rect 414302 161112 414482 161200
rect 426782 161112 426962 161200
rect 427070 161112 427250 161200
rect 427358 161112 427538 161200
rect 427646 161112 427826 161200
rect 427934 161112 428114 161200
rect 428222 161112 428402 161200
rect 428510 161112 428690 161200
rect 428798 161112 428978 161200
rect 441278 161112 441458 161200
rect 441566 161112 441746 161200
rect 441854 161112 442034 161200
rect 442142 161112 442322 161200
rect 442430 161112 442610 161200
rect 442718 161112 442898 161200
rect 443006 161112 443186 161200
rect 443294 161112 443474 161200
rect 455774 161112 455954 161200
rect 456062 161112 456242 161200
rect 456350 161112 456530 161200
rect 456638 161112 456818 161200
rect 456926 161112 457106 161200
rect 457214 161112 457394 161200
rect 457502 161112 457682 161200
rect 457790 161112 457970 161200
rect 180350 160636 180530 160724
rect 180638 160636 180818 160724
rect 180926 160636 181106 160724
rect 181214 160636 181394 160724
rect 181502 160636 181682 160724
rect 181790 160636 181970 160724
rect 182078 160636 182258 160724
rect 182366 160636 182546 160724
rect 194846 160636 195026 160724
rect 195134 160636 195314 160724
rect 195422 160636 195602 160724
rect 195710 160636 195890 160724
rect 195998 160636 196178 160724
rect 196286 160636 196466 160724
rect 196574 160636 196754 160724
rect 196862 160636 197042 160724
rect 209342 160636 209522 160724
rect 209630 160636 209810 160724
rect 209918 160636 210098 160724
rect 210206 160636 210386 160724
rect 210494 160636 210674 160724
rect 210782 160636 210962 160724
rect 211070 160636 211250 160724
rect 211358 160636 211538 160724
rect 223838 160636 224018 160724
rect 224126 160636 224306 160724
rect 224414 160636 224594 160724
rect 224702 160636 224882 160724
rect 224990 160636 225170 160724
rect 225278 160636 225458 160724
rect 225566 160636 225746 160724
rect 225854 160636 226034 160724
rect 238334 160636 238514 160724
rect 238622 160636 238802 160724
rect 238910 160636 239090 160724
rect 239198 160636 239378 160724
rect 239486 160636 239666 160724
rect 239774 160636 239954 160724
rect 240062 160636 240242 160724
rect 240350 160636 240530 160724
rect 252830 160636 253010 160724
rect 253118 160636 253298 160724
rect 253406 160636 253586 160724
rect 253694 160636 253874 160724
rect 253982 160636 254162 160724
rect 254270 160636 254450 160724
rect 254558 160636 254738 160724
rect 254846 160636 255026 160724
rect 267326 160636 267506 160724
rect 267614 160636 267794 160724
rect 267902 160636 268082 160724
rect 268190 160636 268370 160724
rect 268478 160636 268658 160724
rect 268766 160636 268946 160724
rect 269054 160636 269234 160724
rect 269342 160636 269522 160724
rect 281822 160636 282002 160724
rect 282110 160636 282290 160724
rect 282398 160636 282578 160724
rect 282686 160636 282866 160724
rect 282974 160636 283154 160724
rect 283262 160636 283442 160724
rect 283550 160636 283730 160724
rect 283838 160636 284018 160724
rect 296318 160636 296498 160724
rect 296606 160636 296786 160724
rect 296894 160636 297074 160724
rect 297182 160636 297362 160724
rect 297470 160636 297650 160724
rect 297758 160636 297938 160724
rect 298046 160636 298226 160724
rect 298334 160636 298514 160724
rect 310814 160636 310994 160724
rect 311102 160636 311282 160724
rect 311390 160636 311570 160724
rect 311678 160636 311858 160724
rect 311966 160636 312146 160724
rect 312254 160636 312434 160724
rect 312542 160636 312722 160724
rect 312830 160636 313010 160724
rect 325310 160636 325490 160724
rect 325598 160636 325778 160724
rect 325886 160636 326066 160724
rect 326174 160636 326354 160724
rect 326462 160636 326642 160724
rect 326750 160636 326930 160724
rect 327038 160636 327218 160724
rect 327326 160636 327506 160724
rect 339806 160636 339986 160724
rect 340094 160636 340274 160724
rect 340382 160636 340562 160724
rect 340670 160636 340850 160724
rect 340958 160636 341138 160724
rect 341246 160636 341426 160724
rect 341534 160636 341714 160724
rect 341822 160636 342002 160724
rect 354302 160636 354482 160724
rect 354590 160636 354770 160724
rect 354878 160636 355058 160724
rect 355166 160636 355346 160724
rect 355454 160636 355634 160724
rect 355742 160636 355922 160724
rect 356030 160636 356210 160724
rect 356318 160636 356498 160724
rect 368798 160636 368978 160724
rect 369086 160636 369266 160724
rect 369374 160636 369554 160724
rect 369662 160636 369842 160724
rect 369950 160636 370130 160724
rect 370238 160636 370418 160724
rect 370526 160636 370706 160724
rect 370814 160636 370994 160724
rect 383294 160636 383474 160724
rect 383582 160636 383762 160724
rect 383870 160636 384050 160724
rect 384158 160636 384338 160724
rect 384446 160636 384626 160724
rect 384734 160636 384914 160724
rect 385022 160636 385202 160724
rect 385310 160636 385490 160724
rect 397790 160636 397970 160724
rect 398078 160636 398258 160724
rect 398366 160636 398546 160724
rect 398654 160636 398834 160724
rect 398942 160636 399122 160724
rect 399230 160636 399410 160724
rect 399518 160636 399698 160724
rect 399806 160636 399986 160724
rect 412286 160636 412466 160724
rect 412574 160636 412754 160724
rect 412862 160636 413042 160724
rect 413150 160636 413330 160724
rect 413438 160636 413618 160724
rect 413726 160636 413906 160724
rect 414014 160636 414194 160724
rect 414302 160636 414482 160724
rect 426782 160636 426962 160724
rect 427070 160636 427250 160724
rect 427358 160636 427538 160724
rect 427646 160636 427826 160724
rect 427934 160636 428114 160724
rect 428222 160636 428402 160724
rect 428510 160636 428690 160724
rect 428798 160636 428978 160724
rect 441278 160636 441458 160724
rect 441566 160636 441746 160724
rect 441854 160636 442034 160724
rect 442142 160636 442322 160724
rect 442430 160636 442610 160724
rect 442718 160636 442898 160724
rect 443006 160636 443186 160724
rect 443294 160636 443474 160724
rect 455774 160636 455954 160724
rect 456062 160636 456242 160724
rect 456350 160636 456530 160724
rect 456638 160636 456818 160724
rect 456926 160636 457106 160724
rect 457214 160636 457394 160724
rect 457502 160636 457682 160724
rect 457790 160636 457970 160724
rect 180350 160420 180530 160508
rect 180638 160420 180818 160508
rect 180926 160420 181106 160508
rect 181214 160420 181394 160508
rect 181502 160420 181682 160508
rect 181790 160420 181970 160508
rect 182078 160420 182258 160508
rect 182366 160420 182546 160508
rect 194846 160420 195026 160508
rect 195134 160420 195314 160508
rect 195422 160420 195602 160508
rect 195710 160420 195890 160508
rect 195998 160420 196178 160508
rect 196286 160420 196466 160508
rect 196574 160420 196754 160508
rect 196862 160420 197042 160508
rect 209342 160420 209522 160508
rect 209630 160420 209810 160508
rect 209918 160420 210098 160508
rect 210206 160420 210386 160508
rect 210494 160420 210674 160508
rect 210782 160420 210962 160508
rect 211070 160420 211250 160508
rect 211358 160420 211538 160508
rect 223838 160420 224018 160508
rect 224126 160420 224306 160508
rect 224414 160420 224594 160508
rect 224702 160420 224882 160508
rect 224990 160420 225170 160508
rect 225278 160420 225458 160508
rect 225566 160420 225746 160508
rect 225854 160420 226034 160508
rect 238334 160420 238514 160508
rect 238622 160420 238802 160508
rect 238910 160420 239090 160508
rect 239198 160420 239378 160508
rect 239486 160420 239666 160508
rect 239774 160420 239954 160508
rect 240062 160420 240242 160508
rect 240350 160420 240530 160508
rect 252830 160420 253010 160508
rect 253118 160420 253298 160508
rect 253406 160420 253586 160508
rect 253694 160420 253874 160508
rect 253982 160420 254162 160508
rect 254270 160420 254450 160508
rect 254558 160420 254738 160508
rect 254846 160420 255026 160508
rect 267326 160420 267506 160508
rect 267614 160420 267794 160508
rect 267902 160420 268082 160508
rect 268190 160420 268370 160508
rect 268478 160420 268658 160508
rect 268766 160420 268946 160508
rect 269054 160420 269234 160508
rect 269342 160420 269522 160508
rect 281822 160420 282002 160508
rect 282110 160420 282290 160508
rect 282398 160420 282578 160508
rect 282686 160420 282866 160508
rect 282974 160420 283154 160508
rect 283262 160420 283442 160508
rect 283550 160420 283730 160508
rect 283838 160420 284018 160508
rect 296318 160420 296498 160508
rect 296606 160420 296786 160508
rect 296894 160420 297074 160508
rect 297182 160420 297362 160508
rect 297470 160420 297650 160508
rect 297758 160420 297938 160508
rect 298046 160420 298226 160508
rect 298334 160420 298514 160508
rect 310814 160420 310994 160508
rect 311102 160420 311282 160508
rect 311390 160420 311570 160508
rect 311678 160420 311858 160508
rect 311966 160420 312146 160508
rect 312254 160420 312434 160508
rect 312542 160420 312722 160508
rect 312830 160420 313010 160508
rect 325310 160420 325490 160508
rect 325598 160420 325778 160508
rect 325886 160420 326066 160508
rect 326174 160420 326354 160508
rect 326462 160420 326642 160508
rect 326750 160420 326930 160508
rect 327038 160420 327218 160508
rect 327326 160420 327506 160508
rect 339806 160420 339986 160508
rect 340094 160420 340274 160508
rect 340382 160420 340562 160508
rect 340670 160420 340850 160508
rect 340958 160420 341138 160508
rect 341246 160420 341426 160508
rect 341534 160420 341714 160508
rect 341822 160420 342002 160508
rect 354302 160420 354482 160508
rect 354590 160420 354770 160508
rect 354878 160420 355058 160508
rect 355166 160420 355346 160508
rect 355454 160420 355634 160508
rect 355742 160420 355922 160508
rect 356030 160420 356210 160508
rect 356318 160420 356498 160508
rect 368798 160420 368978 160508
rect 369086 160420 369266 160508
rect 369374 160420 369554 160508
rect 369662 160420 369842 160508
rect 369950 160420 370130 160508
rect 370238 160420 370418 160508
rect 370526 160420 370706 160508
rect 370814 160420 370994 160508
rect 383294 160420 383474 160508
rect 383582 160420 383762 160508
rect 383870 160420 384050 160508
rect 384158 160420 384338 160508
rect 384446 160420 384626 160508
rect 384734 160420 384914 160508
rect 385022 160420 385202 160508
rect 385310 160420 385490 160508
rect 397790 160420 397970 160508
rect 398078 160420 398258 160508
rect 398366 160420 398546 160508
rect 398654 160420 398834 160508
rect 398942 160420 399122 160508
rect 399230 160420 399410 160508
rect 399518 160420 399698 160508
rect 399806 160420 399986 160508
rect 412286 160420 412466 160508
rect 412574 160420 412754 160508
rect 412862 160420 413042 160508
rect 413150 160420 413330 160508
rect 413438 160420 413618 160508
rect 413726 160420 413906 160508
rect 414014 160420 414194 160508
rect 414302 160420 414482 160508
rect 426782 160420 426962 160508
rect 427070 160420 427250 160508
rect 427358 160420 427538 160508
rect 427646 160420 427826 160508
rect 427934 160420 428114 160508
rect 428222 160420 428402 160508
rect 428510 160420 428690 160508
rect 428798 160420 428978 160508
rect 441278 160420 441458 160508
rect 441566 160420 441746 160508
rect 441854 160420 442034 160508
rect 442142 160420 442322 160508
rect 442430 160420 442610 160508
rect 442718 160420 442898 160508
rect 443006 160420 443186 160508
rect 443294 160420 443474 160508
rect 455774 160420 455954 160508
rect 456062 160420 456242 160508
rect 456350 160420 456530 160508
rect 456638 160420 456818 160508
rect 456926 160420 457106 160508
rect 457214 160420 457394 160508
rect 457502 160420 457682 160508
rect 457790 160420 457970 160508
rect 180350 146268 180530 146356
rect 180638 146268 180818 146356
rect 180926 146268 181106 146356
rect 181214 146268 181394 146356
rect 181502 146268 181682 146356
rect 181790 146268 181970 146356
rect 182078 146268 182258 146356
rect 182366 146268 182546 146356
rect 194846 146268 195026 146356
rect 195134 146268 195314 146356
rect 195422 146268 195602 146356
rect 195710 146268 195890 146356
rect 195998 146268 196178 146356
rect 196286 146268 196466 146356
rect 196574 146268 196754 146356
rect 196862 146268 197042 146356
rect 209342 146268 209522 146356
rect 209630 146268 209810 146356
rect 209918 146268 210098 146356
rect 210206 146268 210386 146356
rect 210494 146268 210674 146356
rect 210782 146268 210962 146356
rect 211070 146268 211250 146356
rect 211358 146268 211538 146356
rect 223838 146268 224018 146356
rect 224126 146268 224306 146356
rect 224414 146268 224594 146356
rect 224702 146268 224882 146356
rect 224990 146268 225170 146356
rect 225278 146268 225458 146356
rect 225566 146268 225746 146356
rect 225854 146268 226034 146356
rect 238334 146268 238514 146356
rect 238622 146268 238802 146356
rect 238910 146268 239090 146356
rect 239198 146268 239378 146356
rect 239486 146268 239666 146356
rect 239774 146268 239954 146356
rect 240062 146268 240242 146356
rect 240350 146268 240530 146356
rect 252830 146268 253010 146356
rect 253118 146268 253298 146356
rect 253406 146268 253586 146356
rect 253694 146268 253874 146356
rect 253982 146268 254162 146356
rect 254270 146268 254450 146356
rect 254558 146268 254738 146356
rect 254846 146268 255026 146356
rect 267326 146268 267506 146356
rect 267614 146268 267794 146356
rect 267902 146268 268082 146356
rect 268190 146268 268370 146356
rect 268478 146268 268658 146356
rect 268766 146268 268946 146356
rect 269054 146268 269234 146356
rect 269342 146268 269522 146356
rect 281822 146268 282002 146356
rect 282110 146268 282290 146356
rect 282398 146268 282578 146356
rect 282686 146268 282866 146356
rect 282974 146268 283154 146356
rect 283262 146268 283442 146356
rect 283550 146268 283730 146356
rect 283838 146268 284018 146356
rect 296318 146268 296498 146356
rect 296606 146268 296786 146356
rect 296894 146268 297074 146356
rect 297182 146268 297362 146356
rect 297470 146268 297650 146356
rect 297758 146268 297938 146356
rect 298046 146268 298226 146356
rect 298334 146268 298514 146356
rect 310814 146268 310994 146356
rect 311102 146268 311282 146356
rect 311390 146268 311570 146356
rect 311678 146268 311858 146356
rect 311966 146268 312146 146356
rect 312254 146268 312434 146356
rect 312542 146268 312722 146356
rect 312830 146268 313010 146356
rect 325310 146268 325490 146356
rect 325598 146268 325778 146356
rect 325886 146268 326066 146356
rect 326174 146268 326354 146356
rect 326462 146268 326642 146356
rect 326750 146268 326930 146356
rect 327038 146268 327218 146356
rect 327326 146268 327506 146356
rect 339806 146268 339986 146356
rect 340094 146268 340274 146356
rect 340382 146268 340562 146356
rect 340670 146268 340850 146356
rect 340958 146268 341138 146356
rect 341246 146268 341426 146356
rect 341534 146268 341714 146356
rect 341822 146268 342002 146356
rect 354302 146268 354482 146356
rect 354590 146268 354770 146356
rect 354878 146268 355058 146356
rect 355166 146268 355346 146356
rect 355454 146268 355634 146356
rect 355742 146268 355922 146356
rect 356030 146268 356210 146356
rect 356318 146268 356498 146356
rect 368798 146268 368978 146356
rect 369086 146268 369266 146356
rect 369374 146268 369554 146356
rect 369662 146268 369842 146356
rect 369950 146268 370130 146356
rect 370238 146268 370418 146356
rect 370526 146268 370706 146356
rect 370814 146268 370994 146356
rect 383294 146268 383474 146356
rect 383582 146268 383762 146356
rect 383870 146268 384050 146356
rect 384158 146268 384338 146356
rect 384446 146268 384626 146356
rect 384734 146268 384914 146356
rect 385022 146268 385202 146356
rect 385310 146268 385490 146356
rect 397790 146268 397970 146356
rect 398078 146268 398258 146356
rect 398366 146268 398546 146356
rect 398654 146268 398834 146356
rect 398942 146268 399122 146356
rect 399230 146268 399410 146356
rect 399518 146268 399698 146356
rect 399806 146268 399986 146356
rect 412286 146268 412466 146356
rect 412574 146268 412754 146356
rect 412862 146268 413042 146356
rect 413150 146268 413330 146356
rect 413438 146268 413618 146356
rect 413726 146268 413906 146356
rect 414014 146268 414194 146356
rect 414302 146268 414482 146356
rect 426782 146268 426962 146356
rect 427070 146268 427250 146356
rect 427358 146268 427538 146356
rect 427646 146268 427826 146356
rect 427934 146268 428114 146356
rect 428222 146268 428402 146356
rect 428510 146268 428690 146356
rect 428798 146268 428978 146356
rect 441278 146268 441458 146356
rect 441566 146268 441746 146356
rect 441854 146268 442034 146356
rect 442142 146268 442322 146356
rect 442430 146268 442610 146356
rect 442718 146268 442898 146356
rect 443006 146268 443186 146356
rect 443294 146268 443474 146356
rect 455774 146268 455954 146356
rect 456062 146268 456242 146356
rect 456350 146268 456530 146356
rect 456638 146268 456818 146356
rect 456926 146268 457106 146356
rect 457214 146268 457394 146356
rect 457502 146268 457682 146356
rect 457790 146268 457970 146356
rect 180350 146052 180530 146140
rect 180638 146052 180818 146140
rect 180926 146052 181106 146140
rect 181214 146052 181394 146140
rect 181502 146052 181682 146140
rect 181790 146052 181970 146140
rect 182078 146052 182258 146140
rect 182366 146052 182546 146140
rect 194846 146052 195026 146140
rect 195134 146052 195314 146140
rect 195422 146052 195602 146140
rect 195710 146052 195890 146140
rect 195998 146052 196178 146140
rect 196286 146052 196466 146140
rect 196574 146052 196754 146140
rect 196862 146052 197042 146140
rect 209342 146052 209522 146140
rect 209630 146052 209810 146140
rect 209918 146052 210098 146140
rect 210206 146052 210386 146140
rect 210494 146052 210674 146140
rect 210782 146052 210962 146140
rect 211070 146052 211250 146140
rect 211358 146052 211538 146140
rect 223838 146052 224018 146140
rect 224126 146052 224306 146140
rect 224414 146052 224594 146140
rect 224702 146052 224882 146140
rect 224990 146052 225170 146140
rect 225278 146052 225458 146140
rect 225566 146052 225746 146140
rect 225854 146052 226034 146140
rect 238334 146052 238514 146140
rect 238622 146052 238802 146140
rect 238910 146052 239090 146140
rect 239198 146052 239378 146140
rect 239486 146052 239666 146140
rect 239774 146052 239954 146140
rect 240062 146052 240242 146140
rect 240350 146052 240530 146140
rect 252830 146052 253010 146140
rect 253118 146052 253298 146140
rect 253406 146052 253586 146140
rect 253694 146052 253874 146140
rect 253982 146052 254162 146140
rect 254270 146052 254450 146140
rect 254558 146052 254738 146140
rect 254846 146052 255026 146140
rect 267326 146052 267506 146140
rect 267614 146052 267794 146140
rect 267902 146052 268082 146140
rect 268190 146052 268370 146140
rect 268478 146052 268658 146140
rect 268766 146052 268946 146140
rect 269054 146052 269234 146140
rect 269342 146052 269522 146140
rect 281822 146052 282002 146140
rect 282110 146052 282290 146140
rect 282398 146052 282578 146140
rect 282686 146052 282866 146140
rect 282974 146052 283154 146140
rect 283262 146052 283442 146140
rect 283550 146052 283730 146140
rect 283838 146052 284018 146140
rect 296318 146052 296498 146140
rect 296606 146052 296786 146140
rect 296894 146052 297074 146140
rect 297182 146052 297362 146140
rect 297470 146052 297650 146140
rect 297758 146052 297938 146140
rect 298046 146052 298226 146140
rect 298334 146052 298514 146140
rect 310814 146052 310994 146140
rect 311102 146052 311282 146140
rect 311390 146052 311570 146140
rect 311678 146052 311858 146140
rect 311966 146052 312146 146140
rect 312254 146052 312434 146140
rect 312542 146052 312722 146140
rect 312830 146052 313010 146140
rect 325310 146052 325490 146140
rect 325598 146052 325778 146140
rect 325886 146052 326066 146140
rect 326174 146052 326354 146140
rect 326462 146052 326642 146140
rect 326750 146052 326930 146140
rect 327038 146052 327218 146140
rect 327326 146052 327506 146140
rect 339806 146052 339986 146140
rect 340094 146052 340274 146140
rect 340382 146052 340562 146140
rect 340670 146052 340850 146140
rect 340958 146052 341138 146140
rect 341246 146052 341426 146140
rect 341534 146052 341714 146140
rect 341822 146052 342002 146140
rect 354302 146052 354482 146140
rect 354590 146052 354770 146140
rect 354878 146052 355058 146140
rect 355166 146052 355346 146140
rect 355454 146052 355634 146140
rect 355742 146052 355922 146140
rect 356030 146052 356210 146140
rect 356318 146052 356498 146140
rect 368798 146052 368978 146140
rect 369086 146052 369266 146140
rect 369374 146052 369554 146140
rect 369662 146052 369842 146140
rect 369950 146052 370130 146140
rect 370238 146052 370418 146140
rect 370526 146052 370706 146140
rect 370814 146052 370994 146140
rect 383294 146052 383474 146140
rect 383582 146052 383762 146140
rect 383870 146052 384050 146140
rect 384158 146052 384338 146140
rect 384446 146052 384626 146140
rect 384734 146052 384914 146140
rect 385022 146052 385202 146140
rect 385310 146052 385490 146140
rect 397790 146052 397970 146140
rect 398078 146052 398258 146140
rect 398366 146052 398546 146140
rect 398654 146052 398834 146140
rect 398942 146052 399122 146140
rect 399230 146052 399410 146140
rect 399518 146052 399698 146140
rect 399806 146052 399986 146140
rect 412286 146052 412466 146140
rect 412574 146052 412754 146140
rect 412862 146052 413042 146140
rect 413150 146052 413330 146140
rect 413438 146052 413618 146140
rect 413726 146052 413906 146140
rect 414014 146052 414194 146140
rect 414302 146052 414482 146140
rect 426782 146052 426962 146140
rect 427070 146052 427250 146140
rect 427358 146052 427538 146140
rect 427646 146052 427826 146140
rect 427934 146052 428114 146140
rect 428222 146052 428402 146140
rect 428510 146052 428690 146140
rect 428798 146052 428978 146140
rect 441278 146052 441458 146140
rect 441566 146052 441746 146140
rect 441854 146052 442034 146140
rect 442142 146052 442322 146140
rect 442430 146052 442610 146140
rect 442718 146052 442898 146140
rect 443006 146052 443186 146140
rect 443294 146052 443474 146140
rect 455774 146052 455954 146140
rect 456062 146052 456242 146140
rect 456350 146052 456530 146140
rect 456638 146052 456818 146140
rect 456926 146052 457106 146140
rect 457214 146052 457394 146140
rect 457502 146052 457682 146140
rect 457790 146052 457970 146140
rect 180350 145576 180530 145664
rect 180638 145576 180818 145664
rect 180926 145576 181106 145664
rect 181214 145576 181394 145664
rect 181502 145576 181682 145664
rect 181790 145576 181970 145664
rect 182078 145576 182258 145664
rect 182366 145576 182546 145664
rect 194846 145576 195026 145664
rect 195134 145576 195314 145664
rect 195422 145576 195602 145664
rect 195710 145576 195890 145664
rect 195998 145576 196178 145664
rect 196286 145576 196466 145664
rect 196574 145576 196754 145664
rect 196862 145576 197042 145664
rect 209342 145576 209522 145664
rect 209630 145576 209810 145664
rect 209918 145576 210098 145664
rect 210206 145576 210386 145664
rect 210494 145576 210674 145664
rect 210782 145576 210962 145664
rect 211070 145576 211250 145664
rect 211358 145576 211538 145664
rect 223838 145576 224018 145664
rect 224126 145576 224306 145664
rect 224414 145576 224594 145664
rect 224702 145576 224882 145664
rect 224990 145576 225170 145664
rect 225278 145576 225458 145664
rect 225566 145576 225746 145664
rect 225854 145576 226034 145664
rect 238334 145576 238514 145664
rect 238622 145576 238802 145664
rect 238910 145576 239090 145664
rect 239198 145576 239378 145664
rect 239486 145576 239666 145664
rect 239774 145576 239954 145664
rect 240062 145576 240242 145664
rect 240350 145576 240530 145664
rect 252830 145576 253010 145664
rect 253118 145576 253298 145664
rect 253406 145576 253586 145664
rect 253694 145576 253874 145664
rect 253982 145576 254162 145664
rect 254270 145576 254450 145664
rect 254558 145576 254738 145664
rect 254846 145576 255026 145664
rect 267326 145576 267506 145664
rect 267614 145576 267794 145664
rect 267902 145576 268082 145664
rect 268190 145576 268370 145664
rect 268478 145576 268658 145664
rect 268766 145576 268946 145664
rect 269054 145576 269234 145664
rect 269342 145576 269522 145664
rect 281822 145576 282002 145664
rect 282110 145576 282290 145664
rect 282398 145576 282578 145664
rect 282686 145576 282866 145664
rect 282974 145576 283154 145664
rect 283262 145576 283442 145664
rect 283550 145576 283730 145664
rect 283838 145576 284018 145664
rect 296318 145576 296498 145664
rect 296606 145576 296786 145664
rect 296894 145576 297074 145664
rect 297182 145576 297362 145664
rect 297470 145576 297650 145664
rect 297758 145576 297938 145664
rect 298046 145576 298226 145664
rect 298334 145576 298514 145664
rect 310814 145576 310994 145664
rect 311102 145576 311282 145664
rect 311390 145576 311570 145664
rect 311678 145576 311858 145664
rect 311966 145576 312146 145664
rect 312254 145576 312434 145664
rect 312542 145576 312722 145664
rect 312830 145576 313010 145664
rect 325310 145576 325490 145664
rect 325598 145576 325778 145664
rect 325886 145576 326066 145664
rect 326174 145576 326354 145664
rect 326462 145576 326642 145664
rect 326750 145576 326930 145664
rect 327038 145576 327218 145664
rect 327326 145576 327506 145664
rect 339806 145576 339986 145664
rect 340094 145576 340274 145664
rect 340382 145576 340562 145664
rect 340670 145576 340850 145664
rect 340958 145576 341138 145664
rect 341246 145576 341426 145664
rect 341534 145576 341714 145664
rect 341822 145576 342002 145664
rect 354302 145576 354482 145664
rect 354590 145576 354770 145664
rect 354878 145576 355058 145664
rect 355166 145576 355346 145664
rect 355454 145576 355634 145664
rect 355742 145576 355922 145664
rect 356030 145576 356210 145664
rect 356318 145576 356498 145664
rect 368798 145576 368978 145664
rect 369086 145576 369266 145664
rect 369374 145576 369554 145664
rect 369662 145576 369842 145664
rect 369950 145576 370130 145664
rect 370238 145576 370418 145664
rect 370526 145576 370706 145664
rect 370814 145576 370994 145664
rect 383294 145576 383474 145664
rect 383582 145576 383762 145664
rect 383870 145576 384050 145664
rect 384158 145576 384338 145664
rect 384446 145576 384626 145664
rect 384734 145576 384914 145664
rect 385022 145576 385202 145664
rect 385310 145576 385490 145664
rect 397790 145576 397970 145664
rect 398078 145576 398258 145664
rect 398366 145576 398546 145664
rect 398654 145576 398834 145664
rect 398942 145576 399122 145664
rect 399230 145576 399410 145664
rect 399518 145576 399698 145664
rect 399806 145576 399986 145664
rect 412286 145576 412466 145664
rect 412574 145576 412754 145664
rect 412862 145576 413042 145664
rect 413150 145576 413330 145664
rect 413438 145576 413618 145664
rect 413726 145576 413906 145664
rect 414014 145576 414194 145664
rect 414302 145576 414482 145664
rect 426782 145576 426962 145664
rect 427070 145576 427250 145664
rect 427358 145576 427538 145664
rect 427646 145576 427826 145664
rect 427934 145576 428114 145664
rect 428222 145576 428402 145664
rect 428510 145576 428690 145664
rect 428798 145576 428978 145664
rect 441278 145576 441458 145664
rect 441566 145576 441746 145664
rect 441854 145576 442034 145664
rect 442142 145576 442322 145664
rect 442430 145576 442610 145664
rect 442718 145576 442898 145664
rect 443006 145576 443186 145664
rect 443294 145576 443474 145664
rect 455774 145576 455954 145664
rect 456062 145576 456242 145664
rect 456350 145576 456530 145664
rect 456638 145576 456818 145664
rect 456926 145576 457106 145664
rect 457214 145576 457394 145664
rect 457502 145576 457682 145664
rect 457790 145576 457970 145664
rect 180350 145360 180530 145448
rect 180638 145360 180818 145448
rect 180926 145360 181106 145448
rect 181214 145360 181394 145448
rect 181502 145360 181682 145448
rect 181790 145360 181970 145448
rect 182078 145360 182258 145448
rect 182366 145360 182546 145448
rect 194846 145360 195026 145448
rect 195134 145360 195314 145448
rect 195422 145360 195602 145448
rect 195710 145360 195890 145448
rect 195998 145360 196178 145448
rect 196286 145360 196466 145448
rect 196574 145360 196754 145448
rect 196862 145360 197042 145448
rect 209342 145360 209522 145448
rect 209630 145360 209810 145448
rect 209918 145360 210098 145448
rect 210206 145360 210386 145448
rect 210494 145360 210674 145448
rect 210782 145360 210962 145448
rect 211070 145360 211250 145448
rect 211358 145360 211538 145448
rect 223838 145360 224018 145448
rect 224126 145360 224306 145448
rect 224414 145360 224594 145448
rect 224702 145360 224882 145448
rect 224990 145360 225170 145448
rect 225278 145360 225458 145448
rect 225566 145360 225746 145448
rect 225854 145360 226034 145448
rect 238334 145360 238514 145448
rect 238622 145360 238802 145448
rect 238910 145360 239090 145448
rect 239198 145360 239378 145448
rect 239486 145360 239666 145448
rect 239774 145360 239954 145448
rect 240062 145360 240242 145448
rect 240350 145360 240530 145448
rect 252830 145360 253010 145448
rect 253118 145360 253298 145448
rect 253406 145360 253586 145448
rect 253694 145360 253874 145448
rect 253982 145360 254162 145448
rect 254270 145360 254450 145448
rect 254558 145360 254738 145448
rect 254846 145360 255026 145448
rect 267326 145360 267506 145448
rect 267614 145360 267794 145448
rect 267902 145360 268082 145448
rect 268190 145360 268370 145448
rect 268478 145360 268658 145448
rect 268766 145360 268946 145448
rect 269054 145360 269234 145448
rect 269342 145360 269522 145448
rect 281822 145360 282002 145448
rect 282110 145360 282290 145448
rect 282398 145360 282578 145448
rect 282686 145360 282866 145448
rect 282974 145360 283154 145448
rect 283262 145360 283442 145448
rect 283550 145360 283730 145448
rect 283838 145360 284018 145448
rect 296318 145360 296498 145448
rect 296606 145360 296786 145448
rect 296894 145360 297074 145448
rect 297182 145360 297362 145448
rect 297470 145360 297650 145448
rect 297758 145360 297938 145448
rect 298046 145360 298226 145448
rect 298334 145360 298514 145448
rect 310814 145360 310994 145448
rect 311102 145360 311282 145448
rect 311390 145360 311570 145448
rect 311678 145360 311858 145448
rect 311966 145360 312146 145448
rect 312254 145360 312434 145448
rect 312542 145360 312722 145448
rect 312830 145360 313010 145448
rect 325310 145360 325490 145448
rect 325598 145360 325778 145448
rect 325886 145360 326066 145448
rect 326174 145360 326354 145448
rect 326462 145360 326642 145448
rect 326750 145360 326930 145448
rect 327038 145360 327218 145448
rect 327326 145360 327506 145448
rect 339806 145360 339986 145448
rect 340094 145360 340274 145448
rect 340382 145360 340562 145448
rect 340670 145360 340850 145448
rect 340958 145360 341138 145448
rect 341246 145360 341426 145448
rect 341534 145360 341714 145448
rect 341822 145360 342002 145448
rect 354302 145360 354482 145448
rect 354590 145360 354770 145448
rect 354878 145360 355058 145448
rect 355166 145360 355346 145448
rect 355454 145360 355634 145448
rect 355742 145360 355922 145448
rect 356030 145360 356210 145448
rect 356318 145360 356498 145448
rect 368798 145360 368978 145448
rect 369086 145360 369266 145448
rect 369374 145360 369554 145448
rect 369662 145360 369842 145448
rect 369950 145360 370130 145448
rect 370238 145360 370418 145448
rect 370526 145360 370706 145448
rect 370814 145360 370994 145448
rect 383294 145360 383474 145448
rect 383582 145360 383762 145448
rect 383870 145360 384050 145448
rect 384158 145360 384338 145448
rect 384446 145360 384626 145448
rect 384734 145360 384914 145448
rect 385022 145360 385202 145448
rect 385310 145360 385490 145448
rect 397790 145360 397970 145448
rect 398078 145360 398258 145448
rect 398366 145360 398546 145448
rect 398654 145360 398834 145448
rect 398942 145360 399122 145448
rect 399230 145360 399410 145448
rect 399518 145360 399698 145448
rect 399806 145360 399986 145448
rect 412286 145360 412466 145448
rect 412574 145360 412754 145448
rect 412862 145360 413042 145448
rect 413150 145360 413330 145448
rect 413438 145360 413618 145448
rect 413726 145360 413906 145448
rect 414014 145360 414194 145448
rect 414302 145360 414482 145448
rect 426782 145360 426962 145448
rect 427070 145360 427250 145448
rect 427358 145360 427538 145448
rect 427646 145360 427826 145448
rect 427934 145360 428114 145448
rect 428222 145360 428402 145448
rect 428510 145360 428690 145448
rect 428798 145360 428978 145448
rect 441278 145360 441458 145448
rect 441566 145360 441746 145448
rect 441854 145360 442034 145448
rect 442142 145360 442322 145448
rect 442430 145360 442610 145448
rect 442718 145360 442898 145448
rect 443006 145360 443186 145448
rect 443294 145360 443474 145448
rect 455774 145360 455954 145448
rect 456062 145360 456242 145448
rect 456350 145360 456530 145448
rect 456638 145360 456818 145448
rect 456926 145360 457106 145448
rect 457214 145360 457394 145448
rect 457502 145360 457682 145448
rect 457790 145360 457970 145448
rect 180350 131208 180530 131296
rect 180638 131208 180818 131296
rect 180926 131208 181106 131296
rect 181214 131208 181394 131296
rect 181502 131208 181682 131296
rect 181790 131208 181970 131296
rect 182078 131208 182258 131296
rect 182366 131208 182546 131296
rect 194846 131208 195026 131296
rect 195134 131208 195314 131296
rect 195422 131208 195602 131296
rect 195710 131208 195890 131296
rect 195998 131208 196178 131296
rect 196286 131208 196466 131296
rect 196574 131208 196754 131296
rect 196862 131208 197042 131296
rect 209342 131208 209522 131296
rect 209630 131208 209810 131296
rect 209918 131208 210098 131296
rect 210206 131208 210386 131296
rect 210494 131208 210674 131296
rect 210782 131208 210962 131296
rect 211070 131208 211250 131296
rect 211358 131208 211538 131296
rect 223838 131208 224018 131296
rect 224126 131208 224306 131296
rect 224414 131208 224594 131296
rect 224702 131208 224882 131296
rect 224990 131208 225170 131296
rect 225278 131208 225458 131296
rect 225566 131208 225746 131296
rect 225854 131208 226034 131296
rect 238334 131208 238514 131296
rect 238622 131208 238802 131296
rect 238910 131208 239090 131296
rect 239198 131208 239378 131296
rect 239486 131208 239666 131296
rect 239774 131208 239954 131296
rect 240062 131208 240242 131296
rect 240350 131208 240530 131296
rect 252830 131208 253010 131296
rect 253118 131208 253298 131296
rect 253406 131208 253586 131296
rect 253694 131208 253874 131296
rect 253982 131208 254162 131296
rect 254270 131208 254450 131296
rect 254558 131208 254738 131296
rect 254846 131208 255026 131296
rect 267326 131208 267506 131296
rect 267614 131208 267794 131296
rect 267902 131208 268082 131296
rect 268190 131208 268370 131296
rect 268478 131208 268658 131296
rect 268766 131208 268946 131296
rect 269054 131208 269234 131296
rect 269342 131208 269522 131296
rect 281822 131208 282002 131296
rect 282110 131208 282290 131296
rect 282398 131208 282578 131296
rect 282686 131208 282866 131296
rect 282974 131208 283154 131296
rect 283262 131208 283442 131296
rect 283550 131208 283730 131296
rect 283838 131208 284018 131296
rect 296318 131208 296498 131296
rect 296606 131208 296786 131296
rect 296894 131208 297074 131296
rect 297182 131208 297362 131296
rect 297470 131208 297650 131296
rect 297758 131208 297938 131296
rect 298046 131208 298226 131296
rect 298334 131208 298514 131296
rect 310814 131208 310994 131296
rect 311102 131208 311282 131296
rect 311390 131208 311570 131296
rect 311678 131208 311858 131296
rect 311966 131208 312146 131296
rect 312254 131208 312434 131296
rect 312542 131208 312722 131296
rect 312830 131208 313010 131296
rect 325310 131208 325490 131296
rect 325598 131208 325778 131296
rect 325886 131208 326066 131296
rect 326174 131208 326354 131296
rect 326462 131208 326642 131296
rect 326750 131208 326930 131296
rect 327038 131208 327218 131296
rect 327326 131208 327506 131296
rect 339806 131208 339986 131296
rect 340094 131208 340274 131296
rect 340382 131208 340562 131296
rect 340670 131208 340850 131296
rect 340958 131208 341138 131296
rect 341246 131208 341426 131296
rect 341534 131208 341714 131296
rect 341822 131208 342002 131296
rect 354302 131208 354482 131296
rect 354590 131208 354770 131296
rect 354878 131208 355058 131296
rect 355166 131208 355346 131296
rect 355454 131208 355634 131296
rect 355742 131208 355922 131296
rect 356030 131208 356210 131296
rect 356318 131208 356498 131296
rect 368798 131208 368978 131296
rect 369086 131208 369266 131296
rect 369374 131208 369554 131296
rect 369662 131208 369842 131296
rect 369950 131208 370130 131296
rect 370238 131208 370418 131296
rect 370526 131208 370706 131296
rect 370814 131208 370994 131296
rect 383294 131208 383474 131296
rect 383582 131208 383762 131296
rect 383870 131208 384050 131296
rect 384158 131208 384338 131296
rect 384446 131208 384626 131296
rect 384734 131208 384914 131296
rect 385022 131208 385202 131296
rect 385310 131208 385490 131296
rect 397790 131208 397970 131296
rect 398078 131208 398258 131296
rect 398366 131208 398546 131296
rect 398654 131208 398834 131296
rect 398942 131208 399122 131296
rect 399230 131208 399410 131296
rect 399518 131208 399698 131296
rect 399806 131208 399986 131296
rect 412286 131208 412466 131296
rect 412574 131208 412754 131296
rect 412862 131208 413042 131296
rect 413150 131208 413330 131296
rect 413438 131208 413618 131296
rect 413726 131208 413906 131296
rect 414014 131208 414194 131296
rect 414302 131208 414482 131296
rect 426782 131208 426962 131296
rect 427070 131208 427250 131296
rect 427358 131208 427538 131296
rect 427646 131208 427826 131296
rect 427934 131208 428114 131296
rect 428222 131208 428402 131296
rect 428510 131208 428690 131296
rect 428798 131208 428978 131296
rect 441278 131208 441458 131296
rect 441566 131208 441746 131296
rect 441854 131208 442034 131296
rect 442142 131208 442322 131296
rect 442430 131208 442610 131296
rect 442718 131208 442898 131296
rect 443006 131208 443186 131296
rect 443294 131208 443474 131296
rect 455774 131208 455954 131296
rect 456062 131208 456242 131296
rect 456350 131208 456530 131296
rect 456638 131208 456818 131296
rect 456926 131208 457106 131296
rect 457214 131208 457394 131296
rect 457502 131208 457682 131296
rect 457790 131208 457970 131296
rect 180350 130992 180530 131080
rect 180638 130992 180818 131080
rect 180926 130992 181106 131080
rect 181214 130992 181394 131080
rect 181502 130992 181682 131080
rect 181790 130992 181970 131080
rect 182078 130992 182258 131080
rect 182366 130992 182546 131080
rect 194846 130992 195026 131080
rect 195134 130992 195314 131080
rect 195422 130992 195602 131080
rect 195710 130992 195890 131080
rect 195998 130992 196178 131080
rect 196286 130992 196466 131080
rect 196574 130992 196754 131080
rect 196862 130992 197042 131080
rect 209342 130992 209522 131080
rect 209630 130992 209810 131080
rect 209918 130992 210098 131080
rect 210206 130992 210386 131080
rect 210494 130992 210674 131080
rect 210782 130992 210962 131080
rect 211070 130992 211250 131080
rect 211358 130992 211538 131080
rect 223838 130992 224018 131080
rect 224126 130992 224306 131080
rect 224414 130992 224594 131080
rect 224702 130992 224882 131080
rect 224990 130992 225170 131080
rect 225278 130992 225458 131080
rect 225566 130992 225746 131080
rect 225854 130992 226034 131080
rect 238334 130992 238514 131080
rect 238622 130992 238802 131080
rect 238910 130992 239090 131080
rect 239198 130992 239378 131080
rect 239486 130992 239666 131080
rect 239774 130992 239954 131080
rect 240062 130992 240242 131080
rect 240350 130992 240530 131080
rect 252830 130992 253010 131080
rect 253118 130992 253298 131080
rect 253406 130992 253586 131080
rect 253694 130992 253874 131080
rect 253982 130992 254162 131080
rect 254270 130992 254450 131080
rect 254558 130992 254738 131080
rect 254846 130992 255026 131080
rect 267326 130992 267506 131080
rect 267614 130992 267794 131080
rect 267902 130992 268082 131080
rect 268190 130992 268370 131080
rect 268478 130992 268658 131080
rect 268766 130992 268946 131080
rect 269054 130992 269234 131080
rect 269342 130992 269522 131080
rect 281822 130992 282002 131080
rect 282110 130992 282290 131080
rect 282398 130992 282578 131080
rect 282686 130992 282866 131080
rect 282974 130992 283154 131080
rect 283262 130992 283442 131080
rect 283550 130992 283730 131080
rect 283838 130992 284018 131080
rect 296318 130992 296498 131080
rect 296606 130992 296786 131080
rect 296894 130992 297074 131080
rect 297182 130992 297362 131080
rect 297470 130992 297650 131080
rect 297758 130992 297938 131080
rect 298046 130992 298226 131080
rect 298334 130992 298514 131080
rect 310814 130992 310994 131080
rect 311102 130992 311282 131080
rect 311390 130992 311570 131080
rect 311678 130992 311858 131080
rect 311966 130992 312146 131080
rect 312254 130992 312434 131080
rect 312542 130992 312722 131080
rect 312830 130992 313010 131080
rect 325310 130992 325490 131080
rect 325598 130992 325778 131080
rect 325886 130992 326066 131080
rect 326174 130992 326354 131080
rect 326462 130992 326642 131080
rect 326750 130992 326930 131080
rect 327038 130992 327218 131080
rect 327326 130992 327506 131080
rect 339806 130992 339986 131080
rect 340094 130992 340274 131080
rect 340382 130992 340562 131080
rect 340670 130992 340850 131080
rect 340958 130992 341138 131080
rect 341246 130992 341426 131080
rect 341534 130992 341714 131080
rect 341822 130992 342002 131080
rect 354302 130992 354482 131080
rect 354590 130992 354770 131080
rect 354878 130992 355058 131080
rect 355166 130992 355346 131080
rect 355454 130992 355634 131080
rect 355742 130992 355922 131080
rect 356030 130992 356210 131080
rect 356318 130992 356498 131080
rect 368798 130992 368978 131080
rect 369086 130992 369266 131080
rect 369374 130992 369554 131080
rect 369662 130992 369842 131080
rect 369950 130992 370130 131080
rect 370238 130992 370418 131080
rect 370526 130992 370706 131080
rect 370814 130992 370994 131080
rect 383294 130992 383474 131080
rect 383582 130992 383762 131080
rect 383870 130992 384050 131080
rect 384158 130992 384338 131080
rect 384446 130992 384626 131080
rect 384734 130992 384914 131080
rect 385022 130992 385202 131080
rect 385310 130992 385490 131080
rect 397790 130992 397970 131080
rect 398078 130992 398258 131080
rect 398366 130992 398546 131080
rect 398654 130992 398834 131080
rect 398942 130992 399122 131080
rect 399230 130992 399410 131080
rect 399518 130992 399698 131080
rect 399806 130992 399986 131080
rect 412286 130992 412466 131080
rect 412574 130992 412754 131080
rect 412862 130992 413042 131080
rect 413150 130992 413330 131080
rect 413438 130992 413618 131080
rect 413726 130992 413906 131080
rect 414014 130992 414194 131080
rect 414302 130992 414482 131080
rect 426782 130992 426962 131080
rect 427070 130992 427250 131080
rect 427358 130992 427538 131080
rect 427646 130992 427826 131080
rect 427934 130992 428114 131080
rect 428222 130992 428402 131080
rect 428510 130992 428690 131080
rect 428798 130992 428978 131080
rect 441278 130992 441458 131080
rect 441566 130992 441746 131080
rect 441854 130992 442034 131080
rect 442142 130992 442322 131080
rect 442430 130992 442610 131080
rect 442718 130992 442898 131080
rect 443006 130992 443186 131080
rect 443294 130992 443474 131080
rect 455774 130992 455954 131080
rect 456062 130992 456242 131080
rect 456350 130992 456530 131080
rect 456638 130992 456818 131080
rect 456926 130992 457106 131080
rect 457214 130992 457394 131080
rect 457502 130992 457682 131080
rect 457790 130992 457970 131080
rect 180350 130516 180530 130604
rect 180638 130516 180818 130604
rect 180926 130516 181106 130604
rect 181214 130516 181394 130604
rect 181502 130516 181682 130604
rect 181790 130516 181970 130604
rect 182078 130516 182258 130604
rect 182366 130516 182546 130604
rect 194846 130516 195026 130604
rect 195134 130516 195314 130604
rect 195422 130516 195602 130604
rect 195710 130516 195890 130604
rect 195998 130516 196178 130604
rect 196286 130516 196466 130604
rect 196574 130516 196754 130604
rect 196862 130516 197042 130604
rect 209342 130516 209522 130604
rect 209630 130516 209810 130604
rect 209918 130516 210098 130604
rect 210206 130516 210386 130604
rect 210494 130516 210674 130604
rect 210782 130516 210962 130604
rect 211070 130516 211250 130604
rect 211358 130516 211538 130604
rect 223838 130516 224018 130604
rect 224126 130516 224306 130604
rect 224414 130516 224594 130604
rect 224702 130516 224882 130604
rect 224990 130516 225170 130604
rect 225278 130516 225458 130604
rect 225566 130516 225746 130604
rect 225854 130516 226034 130604
rect 238334 130516 238514 130604
rect 238622 130516 238802 130604
rect 238910 130516 239090 130604
rect 239198 130516 239378 130604
rect 239486 130516 239666 130604
rect 239774 130516 239954 130604
rect 240062 130516 240242 130604
rect 240350 130516 240530 130604
rect 252830 130516 253010 130604
rect 253118 130516 253298 130604
rect 253406 130516 253586 130604
rect 253694 130516 253874 130604
rect 253982 130516 254162 130604
rect 254270 130516 254450 130604
rect 254558 130516 254738 130604
rect 254846 130516 255026 130604
rect 267326 130516 267506 130604
rect 267614 130516 267794 130604
rect 267902 130516 268082 130604
rect 268190 130516 268370 130604
rect 268478 130516 268658 130604
rect 268766 130516 268946 130604
rect 269054 130516 269234 130604
rect 269342 130516 269522 130604
rect 281822 130516 282002 130604
rect 282110 130516 282290 130604
rect 282398 130516 282578 130604
rect 282686 130516 282866 130604
rect 282974 130516 283154 130604
rect 283262 130516 283442 130604
rect 283550 130516 283730 130604
rect 283838 130516 284018 130604
rect 296318 130516 296498 130604
rect 296606 130516 296786 130604
rect 296894 130516 297074 130604
rect 297182 130516 297362 130604
rect 297470 130516 297650 130604
rect 297758 130516 297938 130604
rect 298046 130516 298226 130604
rect 298334 130516 298514 130604
rect 310814 130516 310994 130604
rect 311102 130516 311282 130604
rect 311390 130516 311570 130604
rect 311678 130516 311858 130604
rect 311966 130516 312146 130604
rect 312254 130516 312434 130604
rect 312542 130516 312722 130604
rect 312830 130516 313010 130604
rect 325310 130516 325490 130604
rect 325598 130516 325778 130604
rect 325886 130516 326066 130604
rect 326174 130516 326354 130604
rect 326462 130516 326642 130604
rect 326750 130516 326930 130604
rect 327038 130516 327218 130604
rect 327326 130516 327506 130604
rect 339806 130516 339986 130604
rect 340094 130516 340274 130604
rect 340382 130516 340562 130604
rect 340670 130516 340850 130604
rect 340958 130516 341138 130604
rect 341246 130516 341426 130604
rect 341534 130516 341714 130604
rect 341822 130516 342002 130604
rect 354302 130516 354482 130604
rect 354590 130516 354770 130604
rect 354878 130516 355058 130604
rect 355166 130516 355346 130604
rect 355454 130516 355634 130604
rect 355742 130516 355922 130604
rect 356030 130516 356210 130604
rect 356318 130516 356498 130604
rect 368798 130516 368978 130604
rect 369086 130516 369266 130604
rect 369374 130516 369554 130604
rect 369662 130516 369842 130604
rect 369950 130516 370130 130604
rect 370238 130516 370418 130604
rect 370526 130516 370706 130604
rect 370814 130516 370994 130604
rect 383294 130516 383474 130604
rect 383582 130516 383762 130604
rect 383870 130516 384050 130604
rect 384158 130516 384338 130604
rect 384446 130516 384626 130604
rect 384734 130516 384914 130604
rect 385022 130516 385202 130604
rect 385310 130516 385490 130604
rect 397790 130516 397970 130604
rect 398078 130516 398258 130604
rect 398366 130516 398546 130604
rect 398654 130516 398834 130604
rect 398942 130516 399122 130604
rect 399230 130516 399410 130604
rect 399518 130516 399698 130604
rect 399806 130516 399986 130604
rect 412286 130516 412466 130604
rect 412574 130516 412754 130604
rect 412862 130516 413042 130604
rect 413150 130516 413330 130604
rect 413438 130516 413618 130604
rect 413726 130516 413906 130604
rect 414014 130516 414194 130604
rect 414302 130516 414482 130604
rect 426782 130516 426962 130604
rect 427070 130516 427250 130604
rect 427358 130516 427538 130604
rect 427646 130516 427826 130604
rect 427934 130516 428114 130604
rect 428222 130516 428402 130604
rect 428510 130516 428690 130604
rect 428798 130516 428978 130604
rect 441278 130516 441458 130604
rect 441566 130516 441746 130604
rect 441854 130516 442034 130604
rect 442142 130516 442322 130604
rect 442430 130516 442610 130604
rect 442718 130516 442898 130604
rect 443006 130516 443186 130604
rect 443294 130516 443474 130604
rect 455774 130516 455954 130604
rect 456062 130516 456242 130604
rect 456350 130516 456530 130604
rect 456638 130516 456818 130604
rect 456926 130516 457106 130604
rect 457214 130516 457394 130604
rect 457502 130516 457682 130604
rect 457790 130516 457970 130604
rect 180350 130300 180530 130388
rect 180638 130300 180818 130388
rect 180926 130300 181106 130388
rect 181214 130300 181394 130388
rect 181502 130300 181682 130388
rect 181790 130300 181970 130388
rect 182078 130300 182258 130388
rect 182366 130300 182546 130388
rect 194846 130300 195026 130388
rect 195134 130300 195314 130388
rect 195422 130300 195602 130388
rect 195710 130300 195890 130388
rect 195998 130300 196178 130388
rect 196286 130300 196466 130388
rect 196574 130300 196754 130388
rect 196862 130300 197042 130388
rect 209342 130300 209522 130388
rect 209630 130300 209810 130388
rect 209918 130300 210098 130388
rect 210206 130300 210386 130388
rect 210494 130300 210674 130388
rect 210782 130300 210962 130388
rect 211070 130300 211250 130388
rect 211358 130300 211538 130388
rect 223838 130300 224018 130388
rect 224126 130300 224306 130388
rect 224414 130300 224594 130388
rect 224702 130300 224882 130388
rect 224990 130300 225170 130388
rect 225278 130300 225458 130388
rect 225566 130300 225746 130388
rect 225854 130300 226034 130388
rect 238334 130300 238514 130388
rect 238622 130300 238802 130388
rect 238910 130300 239090 130388
rect 239198 130300 239378 130388
rect 239486 130300 239666 130388
rect 239774 130300 239954 130388
rect 240062 130300 240242 130388
rect 240350 130300 240530 130388
rect 252830 130300 253010 130388
rect 253118 130300 253298 130388
rect 253406 130300 253586 130388
rect 253694 130300 253874 130388
rect 253982 130300 254162 130388
rect 254270 130300 254450 130388
rect 254558 130300 254738 130388
rect 254846 130300 255026 130388
rect 267326 130300 267506 130388
rect 267614 130300 267794 130388
rect 267902 130300 268082 130388
rect 268190 130300 268370 130388
rect 268478 130300 268658 130388
rect 268766 130300 268946 130388
rect 269054 130300 269234 130388
rect 269342 130300 269522 130388
rect 281822 130300 282002 130388
rect 282110 130300 282290 130388
rect 282398 130300 282578 130388
rect 282686 130300 282866 130388
rect 282974 130300 283154 130388
rect 283262 130300 283442 130388
rect 283550 130300 283730 130388
rect 283838 130300 284018 130388
rect 296318 130300 296498 130388
rect 296606 130300 296786 130388
rect 296894 130300 297074 130388
rect 297182 130300 297362 130388
rect 297470 130300 297650 130388
rect 297758 130300 297938 130388
rect 298046 130300 298226 130388
rect 298334 130300 298514 130388
rect 310814 130300 310994 130388
rect 311102 130300 311282 130388
rect 311390 130300 311570 130388
rect 311678 130300 311858 130388
rect 311966 130300 312146 130388
rect 312254 130300 312434 130388
rect 312542 130300 312722 130388
rect 312830 130300 313010 130388
rect 325310 130300 325490 130388
rect 325598 130300 325778 130388
rect 325886 130300 326066 130388
rect 326174 130300 326354 130388
rect 326462 130300 326642 130388
rect 326750 130300 326930 130388
rect 327038 130300 327218 130388
rect 327326 130300 327506 130388
rect 339806 130300 339986 130388
rect 340094 130300 340274 130388
rect 340382 130300 340562 130388
rect 340670 130300 340850 130388
rect 340958 130300 341138 130388
rect 341246 130300 341426 130388
rect 341534 130300 341714 130388
rect 341822 130300 342002 130388
rect 354302 130300 354482 130388
rect 354590 130300 354770 130388
rect 354878 130300 355058 130388
rect 355166 130300 355346 130388
rect 355454 130300 355634 130388
rect 355742 130300 355922 130388
rect 356030 130300 356210 130388
rect 356318 130300 356498 130388
rect 368798 130300 368978 130388
rect 369086 130300 369266 130388
rect 369374 130300 369554 130388
rect 369662 130300 369842 130388
rect 369950 130300 370130 130388
rect 370238 130300 370418 130388
rect 370526 130300 370706 130388
rect 370814 130300 370994 130388
rect 383294 130300 383474 130388
rect 383582 130300 383762 130388
rect 383870 130300 384050 130388
rect 384158 130300 384338 130388
rect 384446 130300 384626 130388
rect 384734 130300 384914 130388
rect 385022 130300 385202 130388
rect 385310 130300 385490 130388
rect 397790 130300 397970 130388
rect 398078 130300 398258 130388
rect 398366 130300 398546 130388
rect 398654 130300 398834 130388
rect 398942 130300 399122 130388
rect 399230 130300 399410 130388
rect 399518 130300 399698 130388
rect 399806 130300 399986 130388
rect 412286 130300 412466 130388
rect 412574 130300 412754 130388
rect 412862 130300 413042 130388
rect 413150 130300 413330 130388
rect 413438 130300 413618 130388
rect 413726 130300 413906 130388
rect 414014 130300 414194 130388
rect 414302 130300 414482 130388
rect 426782 130300 426962 130388
rect 427070 130300 427250 130388
rect 427358 130300 427538 130388
rect 427646 130300 427826 130388
rect 427934 130300 428114 130388
rect 428222 130300 428402 130388
rect 428510 130300 428690 130388
rect 428798 130300 428978 130388
rect 441278 130300 441458 130388
rect 441566 130300 441746 130388
rect 441854 130300 442034 130388
rect 442142 130300 442322 130388
rect 442430 130300 442610 130388
rect 442718 130300 442898 130388
rect 443006 130300 443186 130388
rect 443294 130300 443474 130388
rect 455774 130300 455954 130388
rect 456062 130300 456242 130388
rect 456350 130300 456530 130388
rect 456638 130300 456818 130388
rect 456926 130300 457106 130388
rect 457214 130300 457394 130388
rect 457502 130300 457682 130388
rect 457790 130300 457970 130388
rect 180350 116148 180530 116236
rect 180638 116148 180818 116236
rect 180926 116148 181106 116236
rect 181214 116148 181394 116236
rect 181502 116148 181682 116236
rect 181790 116148 181970 116236
rect 182078 116148 182258 116236
rect 182366 116148 182546 116236
rect 194846 116148 195026 116236
rect 195134 116148 195314 116236
rect 195422 116148 195602 116236
rect 195710 116148 195890 116236
rect 195998 116148 196178 116236
rect 196286 116148 196466 116236
rect 196574 116148 196754 116236
rect 196862 116148 197042 116236
rect 209342 116148 209522 116236
rect 209630 116148 209810 116236
rect 209918 116148 210098 116236
rect 210206 116148 210386 116236
rect 210494 116148 210674 116236
rect 210782 116148 210962 116236
rect 211070 116148 211250 116236
rect 211358 116148 211538 116236
rect 223838 116148 224018 116236
rect 224126 116148 224306 116236
rect 224414 116148 224594 116236
rect 224702 116148 224882 116236
rect 224990 116148 225170 116236
rect 225278 116148 225458 116236
rect 225566 116148 225746 116236
rect 225854 116148 226034 116236
rect 238334 116148 238514 116236
rect 238622 116148 238802 116236
rect 238910 116148 239090 116236
rect 239198 116148 239378 116236
rect 239486 116148 239666 116236
rect 239774 116148 239954 116236
rect 240062 116148 240242 116236
rect 240350 116148 240530 116236
rect 252830 116148 253010 116236
rect 253118 116148 253298 116236
rect 253406 116148 253586 116236
rect 253694 116148 253874 116236
rect 253982 116148 254162 116236
rect 254270 116148 254450 116236
rect 254558 116148 254738 116236
rect 254846 116148 255026 116236
rect 267326 116148 267506 116236
rect 267614 116148 267794 116236
rect 267902 116148 268082 116236
rect 268190 116148 268370 116236
rect 268478 116148 268658 116236
rect 268766 116148 268946 116236
rect 269054 116148 269234 116236
rect 269342 116148 269522 116236
rect 281822 116148 282002 116236
rect 282110 116148 282290 116236
rect 282398 116148 282578 116236
rect 282686 116148 282866 116236
rect 282974 116148 283154 116236
rect 283262 116148 283442 116236
rect 283550 116148 283730 116236
rect 283838 116148 284018 116236
rect 296318 116148 296498 116236
rect 296606 116148 296786 116236
rect 296894 116148 297074 116236
rect 297182 116148 297362 116236
rect 297470 116148 297650 116236
rect 297758 116148 297938 116236
rect 298046 116148 298226 116236
rect 298334 116148 298514 116236
rect 310814 116148 310994 116236
rect 311102 116148 311282 116236
rect 311390 116148 311570 116236
rect 311678 116148 311858 116236
rect 311966 116148 312146 116236
rect 312254 116148 312434 116236
rect 312542 116148 312722 116236
rect 312830 116148 313010 116236
rect 325310 116148 325490 116236
rect 325598 116148 325778 116236
rect 325886 116148 326066 116236
rect 326174 116148 326354 116236
rect 326462 116148 326642 116236
rect 326750 116148 326930 116236
rect 327038 116148 327218 116236
rect 327326 116148 327506 116236
rect 339806 116148 339986 116236
rect 340094 116148 340274 116236
rect 340382 116148 340562 116236
rect 340670 116148 340850 116236
rect 340958 116148 341138 116236
rect 341246 116148 341426 116236
rect 341534 116148 341714 116236
rect 341822 116148 342002 116236
rect 354302 116148 354482 116236
rect 354590 116148 354770 116236
rect 354878 116148 355058 116236
rect 355166 116148 355346 116236
rect 355454 116148 355634 116236
rect 355742 116148 355922 116236
rect 356030 116148 356210 116236
rect 356318 116148 356498 116236
rect 368798 116148 368978 116236
rect 369086 116148 369266 116236
rect 369374 116148 369554 116236
rect 369662 116148 369842 116236
rect 369950 116148 370130 116236
rect 370238 116148 370418 116236
rect 370526 116148 370706 116236
rect 370814 116148 370994 116236
rect 383294 116148 383474 116236
rect 383582 116148 383762 116236
rect 383870 116148 384050 116236
rect 384158 116148 384338 116236
rect 384446 116148 384626 116236
rect 384734 116148 384914 116236
rect 385022 116148 385202 116236
rect 385310 116148 385490 116236
rect 397790 116148 397970 116236
rect 398078 116148 398258 116236
rect 398366 116148 398546 116236
rect 398654 116148 398834 116236
rect 398942 116148 399122 116236
rect 399230 116148 399410 116236
rect 399518 116148 399698 116236
rect 399806 116148 399986 116236
rect 412286 116148 412466 116236
rect 412574 116148 412754 116236
rect 412862 116148 413042 116236
rect 413150 116148 413330 116236
rect 413438 116148 413618 116236
rect 413726 116148 413906 116236
rect 414014 116148 414194 116236
rect 414302 116148 414482 116236
rect 426782 116148 426962 116236
rect 427070 116148 427250 116236
rect 427358 116148 427538 116236
rect 427646 116148 427826 116236
rect 427934 116148 428114 116236
rect 428222 116148 428402 116236
rect 428510 116148 428690 116236
rect 428798 116148 428978 116236
rect 441278 116148 441458 116236
rect 441566 116148 441746 116236
rect 441854 116148 442034 116236
rect 442142 116148 442322 116236
rect 442430 116148 442610 116236
rect 442718 116148 442898 116236
rect 443006 116148 443186 116236
rect 443294 116148 443474 116236
rect 455774 116148 455954 116236
rect 456062 116148 456242 116236
rect 456350 116148 456530 116236
rect 456638 116148 456818 116236
rect 456926 116148 457106 116236
rect 457214 116148 457394 116236
rect 457502 116148 457682 116236
rect 457790 116148 457970 116236
rect 180350 115932 180530 116020
rect 180638 115932 180818 116020
rect 180926 115932 181106 116020
rect 181214 115932 181394 116020
rect 181502 115932 181682 116020
rect 181790 115932 181970 116020
rect 182078 115932 182258 116020
rect 182366 115932 182546 116020
rect 194846 115932 195026 116020
rect 195134 115932 195314 116020
rect 195422 115932 195602 116020
rect 195710 115932 195890 116020
rect 195998 115932 196178 116020
rect 196286 115932 196466 116020
rect 196574 115932 196754 116020
rect 196862 115932 197042 116020
rect 209342 115932 209522 116020
rect 209630 115932 209810 116020
rect 209918 115932 210098 116020
rect 210206 115932 210386 116020
rect 210494 115932 210674 116020
rect 210782 115932 210962 116020
rect 211070 115932 211250 116020
rect 211358 115932 211538 116020
rect 223838 115932 224018 116020
rect 224126 115932 224306 116020
rect 224414 115932 224594 116020
rect 224702 115932 224882 116020
rect 224990 115932 225170 116020
rect 225278 115932 225458 116020
rect 225566 115932 225746 116020
rect 225854 115932 226034 116020
rect 238334 115932 238514 116020
rect 238622 115932 238802 116020
rect 238910 115932 239090 116020
rect 239198 115932 239378 116020
rect 239486 115932 239666 116020
rect 239774 115932 239954 116020
rect 240062 115932 240242 116020
rect 240350 115932 240530 116020
rect 252830 115932 253010 116020
rect 253118 115932 253298 116020
rect 253406 115932 253586 116020
rect 253694 115932 253874 116020
rect 253982 115932 254162 116020
rect 254270 115932 254450 116020
rect 254558 115932 254738 116020
rect 254846 115932 255026 116020
rect 267326 115932 267506 116020
rect 267614 115932 267794 116020
rect 267902 115932 268082 116020
rect 268190 115932 268370 116020
rect 268478 115932 268658 116020
rect 268766 115932 268946 116020
rect 269054 115932 269234 116020
rect 269342 115932 269522 116020
rect 281822 115932 282002 116020
rect 282110 115932 282290 116020
rect 282398 115932 282578 116020
rect 282686 115932 282866 116020
rect 282974 115932 283154 116020
rect 283262 115932 283442 116020
rect 283550 115932 283730 116020
rect 283838 115932 284018 116020
rect 296318 115932 296498 116020
rect 296606 115932 296786 116020
rect 296894 115932 297074 116020
rect 297182 115932 297362 116020
rect 297470 115932 297650 116020
rect 297758 115932 297938 116020
rect 298046 115932 298226 116020
rect 298334 115932 298514 116020
rect 310814 115932 310994 116020
rect 311102 115932 311282 116020
rect 311390 115932 311570 116020
rect 311678 115932 311858 116020
rect 311966 115932 312146 116020
rect 312254 115932 312434 116020
rect 312542 115932 312722 116020
rect 312830 115932 313010 116020
rect 325310 115932 325490 116020
rect 325598 115932 325778 116020
rect 325886 115932 326066 116020
rect 326174 115932 326354 116020
rect 326462 115932 326642 116020
rect 326750 115932 326930 116020
rect 327038 115932 327218 116020
rect 327326 115932 327506 116020
rect 339806 115932 339986 116020
rect 340094 115932 340274 116020
rect 340382 115932 340562 116020
rect 340670 115932 340850 116020
rect 340958 115932 341138 116020
rect 341246 115932 341426 116020
rect 341534 115932 341714 116020
rect 341822 115932 342002 116020
rect 354302 115932 354482 116020
rect 354590 115932 354770 116020
rect 354878 115932 355058 116020
rect 355166 115932 355346 116020
rect 355454 115932 355634 116020
rect 355742 115932 355922 116020
rect 356030 115932 356210 116020
rect 356318 115932 356498 116020
rect 368798 115932 368978 116020
rect 369086 115932 369266 116020
rect 369374 115932 369554 116020
rect 369662 115932 369842 116020
rect 369950 115932 370130 116020
rect 370238 115932 370418 116020
rect 370526 115932 370706 116020
rect 370814 115932 370994 116020
rect 383294 115932 383474 116020
rect 383582 115932 383762 116020
rect 383870 115932 384050 116020
rect 384158 115932 384338 116020
rect 384446 115932 384626 116020
rect 384734 115932 384914 116020
rect 385022 115932 385202 116020
rect 385310 115932 385490 116020
rect 397790 115932 397970 116020
rect 398078 115932 398258 116020
rect 398366 115932 398546 116020
rect 398654 115932 398834 116020
rect 398942 115932 399122 116020
rect 399230 115932 399410 116020
rect 399518 115932 399698 116020
rect 399806 115932 399986 116020
rect 412286 115932 412466 116020
rect 412574 115932 412754 116020
rect 412862 115932 413042 116020
rect 413150 115932 413330 116020
rect 413438 115932 413618 116020
rect 413726 115932 413906 116020
rect 414014 115932 414194 116020
rect 414302 115932 414482 116020
rect 426782 115932 426962 116020
rect 427070 115932 427250 116020
rect 427358 115932 427538 116020
rect 427646 115932 427826 116020
rect 427934 115932 428114 116020
rect 428222 115932 428402 116020
rect 428510 115932 428690 116020
rect 428798 115932 428978 116020
rect 441278 115932 441458 116020
rect 441566 115932 441746 116020
rect 441854 115932 442034 116020
rect 442142 115932 442322 116020
rect 442430 115932 442610 116020
rect 442718 115932 442898 116020
rect 443006 115932 443186 116020
rect 443294 115932 443474 116020
rect 455774 115932 455954 116020
rect 456062 115932 456242 116020
rect 456350 115932 456530 116020
rect 456638 115932 456818 116020
rect 456926 115932 457106 116020
rect 457214 115932 457394 116020
rect 457502 115932 457682 116020
rect 457790 115932 457970 116020
rect 180350 115456 180530 115544
rect 180638 115456 180818 115544
rect 180926 115456 181106 115544
rect 181214 115456 181394 115544
rect 181502 115456 181682 115544
rect 181790 115456 181970 115544
rect 182078 115456 182258 115544
rect 182366 115456 182546 115544
rect 194846 115456 195026 115544
rect 195134 115456 195314 115544
rect 195422 115456 195602 115544
rect 195710 115456 195890 115544
rect 195998 115456 196178 115544
rect 196286 115456 196466 115544
rect 196574 115456 196754 115544
rect 196862 115456 197042 115544
rect 209342 115456 209522 115544
rect 209630 115456 209810 115544
rect 209918 115456 210098 115544
rect 210206 115456 210386 115544
rect 210494 115456 210674 115544
rect 210782 115456 210962 115544
rect 211070 115456 211250 115544
rect 211358 115456 211538 115544
rect 223838 115456 224018 115544
rect 224126 115456 224306 115544
rect 224414 115456 224594 115544
rect 224702 115456 224882 115544
rect 224990 115456 225170 115544
rect 225278 115456 225458 115544
rect 225566 115456 225746 115544
rect 225854 115456 226034 115544
rect 238334 115456 238514 115544
rect 238622 115456 238802 115544
rect 238910 115456 239090 115544
rect 239198 115456 239378 115544
rect 239486 115456 239666 115544
rect 239774 115456 239954 115544
rect 240062 115456 240242 115544
rect 240350 115456 240530 115544
rect 252830 115456 253010 115544
rect 253118 115456 253298 115544
rect 253406 115456 253586 115544
rect 253694 115456 253874 115544
rect 253982 115456 254162 115544
rect 254270 115456 254450 115544
rect 254558 115456 254738 115544
rect 254846 115456 255026 115544
rect 267326 115456 267506 115544
rect 267614 115456 267794 115544
rect 267902 115456 268082 115544
rect 268190 115456 268370 115544
rect 268478 115456 268658 115544
rect 268766 115456 268946 115544
rect 269054 115456 269234 115544
rect 269342 115456 269522 115544
rect 281822 115456 282002 115544
rect 282110 115456 282290 115544
rect 282398 115456 282578 115544
rect 282686 115456 282866 115544
rect 282974 115456 283154 115544
rect 283262 115456 283442 115544
rect 283550 115456 283730 115544
rect 283838 115456 284018 115544
rect 296318 115456 296498 115544
rect 296606 115456 296786 115544
rect 296894 115456 297074 115544
rect 297182 115456 297362 115544
rect 297470 115456 297650 115544
rect 297758 115456 297938 115544
rect 298046 115456 298226 115544
rect 298334 115456 298514 115544
rect 310814 115456 310994 115544
rect 311102 115456 311282 115544
rect 311390 115456 311570 115544
rect 311678 115456 311858 115544
rect 311966 115456 312146 115544
rect 312254 115456 312434 115544
rect 312542 115456 312722 115544
rect 312830 115456 313010 115544
rect 325310 115456 325490 115544
rect 325598 115456 325778 115544
rect 325886 115456 326066 115544
rect 326174 115456 326354 115544
rect 326462 115456 326642 115544
rect 326750 115456 326930 115544
rect 327038 115456 327218 115544
rect 327326 115456 327506 115544
rect 339806 115456 339986 115544
rect 340094 115456 340274 115544
rect 340382 115456 340562 115544
rect 340670 115456 340850 115544
rect 340958 115456 341138 115544
rect 341246 115456 341426 115544
rect 341534 115456 341714 115544
rect 341822 115456 342002 115544
rect 354302 115456 354482 115544
rect 354590 115456 354770 115544
rect 354878 115456 355058 115544
rect 355166 115456 355346 115544
rect 355454 115456 355634 115544
rect 355742 115456 355922 115544
rect 356030 115456 356210 115544
rect 356318 115456 356498 115544
rect 368798 115456 368978 115544
rect 369086 115456 369266 115544
rect 369374 115456 369554 115544
rect 369662 115456 369842 115544
rect 369950 115456 370130 115544
rect 370238 115456 370418 115544
rect 370526 115456 370706 115544
rect 370814 115456 370994 115544
rect 383294 115456 383474 115544
rect 383582 115456 383762 115544
rect 383870 115456 384050 115544
rect 384158 115456 384338 115544
rect 384446 115456 384626 115544
rect 384734 115456 384914 115544
rect 385022 115456 385202 115544
rect 385310 115456 385490 115544
rect 397790 115456 397970 115544
rect 398078 115456 398258 115544
rect 398366 115456 398546 115544
rect 398654 115456 398834 115544
rect 398942 115456 399122 115544
rect 399230 115456 399410 115544
rect 399518 115456 399698 115544
rect 399806 115456 399986 115544
rect 412286 115456 412466 115544
rect 412574 115456 412754 115544
rect 412862 115456 413042 115544
rect 413150 115456 413330 115544
rect 413438 115456 413618 115544
rect 413726 115456 413906 115544
rect 414014 115456 414194 115544
rect 414302 115456 414482 115544
rect 426782 115456 426962 115544
rect 427070 115456 427250 115544
rect 427358 115456 427538 115544
rect 427646 115456 427826 115544
rect 427934 115456 428114 115544
rect 428222 115456 428402 115544
rect 428510 115456 428690 115544
rect 428798 115456 428978 115544
rect 441278 115456 441458 115544
rect 441566 115456 441746 115544
rect 441854 115456 442034 115544
rect 442142 115456 442322 115544
rect 442430 115456 442610 115544
rect 442718 115456 442898 115544
rect 443006 115456 443186 115544
rect 443294 115456 443474 115544
rect 455774 115456 455954 115544
rect 456062 115456 456242 115544
rect 456350 115456 456530 115544
rect 456638 115456 456818 115544
rect 456926 115456 457106 115544
rect 457214 115456 457394 115544
rect 457502 115456 457682 115544
rect 457790 115456 457970 115544
rect 180350 115240 180530 115328
rect 180638 115240 180818 115328
rect 180926 115240 181106 115328
rect 181214 115240 181394 115328
rect 181502 115240 181682 115328
rect 181790 115240 181970 115328
rect 182078 115240 182258 115328
rect 182366 115240 182546 115328
rect 194846 115240 195026 115328
rect 195134 115240 195314 115328
rect 195422 115240 195602 115328
rect 195710 115240 195890 115328
rect 195998 115240 196178 115328
rect 196286 115240 196466 115328
rect 196574 115240 196754 115328
rect 196862 115240 197042 115328
rect 209342 115240 209522 115328
rect 209630 115240 209810 115328
rect 209918 115240 210098 115328
rect 210206 115240 210386 115328
rect 210494 115240 210674 115328
rect 210782 115240 210962 115328
rect 211070 115240 211250 115328
rect 211358 115240 211538 115328
rect 223838 115240 224018 115328
rect 224126 115240 224306 115328
rect 224414 115240 224594 115328
rect 224702 115240 224882 115328
rect 224990 115240 225170 115328
rect 225278 115240 225458 115328
rect 225566 115240 225746 115328
rect 225854 115240 226034 115328
rect 238334 115240 238514 115328
rect 238622 115240 238802 115328
rect 238910 115240 239090 115328
rect 239198 115240 239378 115328
rect 239486 115240 239666 115328
rect 239774 115240 239954 115328
rect 240062 115240 240242 115328
rect 240350 115240 240530 115328
rect 252830 115240 253010 115328
rect 253118 115240 253298 115328
rect 253406 115240 253586 115328
rect 253694 115240 253874 115328
rect 253982 115240 254162 115328
rect 254270 115240 254450 115328
rect 254558 115240 254738 115328
rect 254846 115240 255026 115328
rect 267326 115240 267506 115328
rect 267614 115240 267794 115328
rect 267902 115240 268082 115328
rect 268190 115240 268370 115328
rect 268478 115240 268658 115328
rect 268766 115240 268946 115328
rect 269054 115240 269234 115328
rect 269342 115240 269522 115328
rect 281822 115240 282002 115328
rect 282110 115240 282290 115328
rect 282398 115240 282578 115328
rect 282686 115240 282866 115328
rect 282974 115240 283154 115328
rect 283262 115240 283442 115328
rect 283550 115240 283730 115328
rect 283838 115240 284018 115328
rect 296318 115240 296498 115328
rect 296606 115240 296786 115328
rect 296894 115240 297074 115328
rect 297182 115240 297362 115328
rect 297470 115240 297650 115328
rect 297758 115240 297938 115328
rect 298046 115240 298226 115328
rect 298334 115240 298514 115328
rect 310814 115240 310994 115328
rect 311102 115240 311282 115328
rect 311390 115240 311570 115328
rect 311678 115240 311858 115328
rect 311966 115240 312146 115328
rect 312254 115240 312434 115328
rect 312542 115240 312722 115328
rect 312830 115240 313010 115328
rect 325310 115240 325490 115328
rect 325598 115240 325778 115328
rect 325886 115240 326066 115328
rect 326174 115240 326354 115328
rect 326462 115240 326642 115328
rect 326750 115240 326930 115328
rect 327038 115240 327218 115328
rect 327326 115240 327506 115328
rect 339806 115240 339986 115328
rect 340094 115240 340274 115328
rect 340382 115240 340562 115328
rect 340670 115240 340850 115328
rect 340958 115240 341138 115328
rect 341246 115240 341426 115328
rect 341534 115240 341714 115328
rect 341822 115240 342002 115328
rect 354302 115240 354482 115328
rect 354590 115240 354770 115328
rect 354878 115240 355058 115328
rect 355166 115240 355346 115328
rect 355454 115240 355634 115328
rect 355742 115240 355922 115328
rect 356030 115240 356210 115328
rect 356318 115240 356498 115328
rect 368798 115240 368978 115328
rect 369086 115240 369266 115328
rect 369374 115240 369554 115328
rect 369662 115240 369842 115328
rect 369950 115240 370130 115328
rect 370238 115240 370418 115328
rect 370526 115240 370706 115328
rect 370814 115240 370994 115328
rect 383294 115240 383474 115328
rect 383582 115240 383762 115328
rect 383870 115240 384050 115328
rect 384158 115240 384338 115328
rect 384446 115240 384626 115328
rect 384734 115240 384914 115328
rect 385022 115240 385202 115328
rect 385310 115240 385490 115328
rect 397790 115240 397970 115328
rect 398078 115240 398258 115328
rect 398366 115240 398546 115328
rect 398654 115240 398834 115328
rect 398942 115240 399122 115328
rect 399230 115240 399410 115328
rect 399518 115240 399698 115328
rect 399806 115240 399986 115328
rect 412286 115240 412466 115328
rect 412574 115240 412754 115328
rect 412862 115240 413042 115328
rect 413150 115240 413330 115328
rect 413438 115240 413618 115328
rect 413726 115240 413906 115328
rect 414014 115240 414194 115328
rect 414302 115240 414482 115328
rect 426782 115240 426962 115328
rect 427070 115240 427250 115328
rect 427358 115240 427538 115328
rect 427646 115240 427826 115328
rect 427934 115240 428114 115328
rect 428222 115240 428402 115328
rect 428510 115240 428690 115328
rect 428798 115240 428978 115328
rect 441278 115240 441458 115328
rect 441566 115240 441746 115328
rect 441854 115240 442034 115328
rect 442142 115240 442322 115328
rect 442430 115240 442610 115328
rect 442718 115240 442898 115328
rect 443006 115240 443186 115328
rect 443294 115240 443474 115328
rect 455774 115240 455954 115328
rect 456062 115240 456242 115328
rect 456350 115240 456530 115328
rect 456638 115240 456818 115328
rect 456926 115240 457106 115328
rect 457214 115240 457394 115328
rect 457502 115240 457682 115328
rect 457790 115240 457970 115328
rect 180350 101088 180530 101176
rect 180638 101088 180818 101176
rect 180926 101088 181106 101176
rect 181214 101088 181394 101176
rect 181502 101088 181682 101176
rect 181790 101088 181970 101176
rect 182078 101088 182258 101176
rect 182366 101088 182546 101176
rect 194846 101088 195026 101176
rect 195134 101088 195314 101176
rect 195422 101088 195602 101176
rect 195710 101088 195890 101176
rect 195998 101088 196178 101176
rect 196286 101088 196466 101176
rect 196574 101088 196754 101176
rect 196862 101088 197042 101176
rect 209342 101088 209522 101176
rect 209630 101088 209810 101176
rect 209918 101088 210098 101176
rect 210206 101088 210386 101176
rect 210494 101088 210674 101176
rect 210782 101088 210962 101176
rect 211070 101088 211250 101176
rect 211358 101088 211538 101176
rect 223838 101088 224018 101176
rect 224126 101088 224306 101176
rect 224414 101088 224594 101176
rect 224702 101088 224882 101176
rect 224990 101088 225170 101176
rect 225278 101088 225458 101176
rect 225566 101088 225746 101176
rect 225854 101088 226034 101176
rect 238334 101088 238514 101176
rect 238622 101088 238802 101176
rect 238910 101088 239090 101176
rect 239198 101088 239378 101176
rect 239486 101088 239666 101176
rect 239774 101088 239954 101176
rect 240062 101088 240242 101176
rect 240350 101088 240530 101176
rect 252830 101088 253010 101176
rect 253118 101088 253298 101176
rect 253406 101088 253586 101176
rect 253694 101088 253874 101176
rect 253982 101088 254162 101176
rect 254270 101088 254450 101176
rect 254558 101088 254738 101176
rect 254846 101088 255026 101176
rect 267326 101088 267506 101176
rect 267614 101088 267794 101176
rect 267902 101088 268082 101176
rect 268190 101088 268370 101176
rect 268478 101088 268658 101176
rect 268766 101088 268946 101176
rect 269054 101088 269234 101176
rect 269342 101088 269522 101176
rect 281822 101088 282002 101176
rect 282110 101088 282290 101176
rect 282398 101088 282578 101176
rect 282686 101088 282866 101176
rect 282974 101088 283154 101176
rect 283262 101088 283442 101176
rect 283550 101088 283730 101176
rect 283838 101088 284018 101176
rect 296318 101088 296498 101176
rect 296606 101088 296786 101176
rect 296894 101088 297074 101176
rect 297182 101088 297362 101176
rect 297470 101088 297650 101176
rect 297758 101088 297938 101176
rect 298046 101088 298226 101176
rect 298334 101088 298514 101176
rect 310814 101088 310994 101176
rect 311102 101088 311282 101176
rect 311390 101088 311570 101176
rect 311678 101088 311858 101176
rect 311966 101088 312146 101176
rect 312254 101088 312434 101176
rect 312542 101088 312722 101176
rect 312830 101088 313010 101176
rect 325310 101088 325490 101176
rect 325598 101088 325778 101176
rect 325886 101088 326066 101176
rect 326174 101088 326354 101176
rect 326462 101088 326642 101176
rect 326750 101088 326930 101176
rect 327038 101088 327218 101176
rect 327326 101088 327506 101176
rect 339806 101088 339986 101176
rect 340094 101088 340274 101176
rect 340382 101088 340562 101176
rect 340670 101088 340850 101176
rect 340958 101088 341138 101176
rect 341246 101088 341426 101176
rect 341534 101088 341714 101176
rect 341822 101088 342002 101176
rect 354302 101088 354482 101176
rect 354590 101088 354770 101176
rect 354878 101088 355058 101176
rect 355166 101088 355346 101176
rect 355454 101088 355634 101176
rect 355742 101088 355922 101176
rect 356030 101088 356210 101176
rect 356318 101088 356498 101176
rect 368798 101088 368978 101176
rect 369086 101088 369266 101176
rect 369374 101088 369554 101176
rect 369662 101088 369842 101176
rect 369950 101088 370130 101176
rect 370238 101088 370418 101176
rect 370526 101088 370706 101176
rect 370814 101088 370994 101176
rect 383294 101088 383474 101176
rect 383582 101088 383762 101176
rect 383870 101088 384050 101176
rect 384158 101088 384338 101176
rect 384446 101088 384626 101176
rect 384734 101088 384914 101176
rect 385022 101088 385202 101176
rect 385310 101088 385490 101176
rect 397790 101088 397970 101176
rect 398078 101088 398258 101176
rect 398366 101088 398546 101176
rect 398654 101088 398834 101176
rect 398942 101088 399122 101176
rect 399230 101088 399410 101176
rect 399518 101088 399698 101176
rect 399806 101088 399986 101176
rect 412286 101088 412466 101176
rect 412574 101088 412754 101176
rect 412862 101088 413042 101176
rect 413150 101088 413330 101176
rect 413438 101088 413618 101176
rect 413726 101088 413906 101176
rect 414014 101088 414194 101176
rect 414302 101088 414482 101176
rect 426782 101088 426962 101176
rect 427070 101088 427250 101176
rect 427358 101088 427538 101176
rect 427646 101088 427826 101176
rect 427934 101088 428114 101176
rect 428222 101088 428402 101176
rect 428510 101088 428690 101176
rect 428798 101088 428978 101176
rect 441278 101088 441458 101176
rect 441566 101088 441746 101176
rect 441854 101088 442034 101176
rect 442142 101088 442322 101176
rect 442430 101088 442610 101176
rect 442718 101088 442898 101176
rect 443006 101088 443186 101176
rect 443294 101088 443474 101176
rect 455774 101088 455954 101176
rect 456062 101088 456242 101176
rect 456350 101088 456530 101176
rect 456638 101088 456818 101176
rect 456926 101088 457106 101176
rect 457214 101088 457394 101176
rect 457502 101088 457682 101176
rect 457790 101088 457970 101176
rect 180350 100872 180530 100960
rect 180638 100872 180818 100960
rect 180926 100872 181106 100960
rect 181214 100872 181394 100960
rect 181502 100872 181682 100960
rect 181790 100872 181970 100960
rect 182078 100872 182258 100960
rect 182366 100872 182546 100960
rect 194846 100872 195026 100960
rect 195134 100872 195314 100960
rect 195422 100872 195602 100960
rect 195710 100872 195890 100960
rect 195998 100872 196178 100960
rect 196286 100872 196466 100960
rect 196574 100872 196754 100960
rect 196862 100872 197042 100960
rect 209342 100872 209522 100960
rect 209630 100872 209810 100960
rect 209918 100872 210098 100960
rect 210206 100872 210386 100960
rect 210494 100872 210674 100960
rect 210782 100872 210962 100960
rect 211070 100872 211250 100960
rect 211358 100872 211538 100960
rect 223838 100872 224018 100960
rect 224126 100872 224306 100960
rect 224414 100872 224594 100960
rect 224702 100872 224882 100960
rect 224990 100872 225170 100960
rect 225278 100872 225458 100960
rect 225566 100872 225746 100960
rect 225854 100872 226034 100960
rect 238334 100872 238514 100960
rect 238622 100872 238802 100960
rect 238910 100872 239090 100960
rect 239198 100872 239378 100960
rect 239486 100872 239666 100960
rect 239774 100872 239954 100960
rect 240062 100872 240242 100960
rect 240350 100872 240530 100960
rect 252830 100872 253010 100960
rect 253118 100872 253298 100960
rect 253406 100872 253586 100960
rect 253694 100872 253874 100960
rect 253982 100872 254162 100960
rect 254270 100872 254450 100960
rect 254558 100872 254738 100960
rect 254846 100872 255026 100960
rect 267326 100872 267506 100960
rect 267614 100872 267794 100960
rect 267902 100872 268082 100960
rect 268190 100872 268370 100960
rect 268478 100872 268658 100960
rect 268766 100872 268946 100960
rect 269054 100872 269234 100960
rect 269342 100872 269522 100960
rect 281822 100872 282002 100960
rect 282110 100872 282290 100960
rect 282398 100872 282578 100960
rect 282686 100872 282866 100960
rect 282974 100872 283154 100960
rect 283262 100872 283442 100960
rect 283550 100872 283730 100960
rect 283838 100872 284018 100960
rect 296318 100872 296498 100960
rect 296606 100872 296786 100960
rect 296894 100872 297074 100960
rect 297182 100872 297362 100960
rect 297470 100872 297650 100960
rect 297758 100872 297938 100960
rect 298046 100872 298226 100960
rect 298334 100872 298514 100960
rect 310814 100872 310994 100960
rect 311102 100872 311282 100960
rect 311390 100872 311570 100960
rect 311678 100872 311858 100960
rect 311966 100872 312146 100960
rect 312254 100872 312434 100960
rect 312542 100872 312722 100960
rect 312830 100872 313010 100960
rect 325310 100872 325490 100960
rect 325598 100872 325778 100960
rect 325886 100872 326066 100960
rect 326174 100872 326354 100960
rect 326462 100872 326642 100960
rect 326750 100872 326930 100960
rect 327038 100872 327218 100960
rect 327326 100872 327506 100960
rect 339806 100872 339986 100960
rect 340094 100872 340274 100960
rect 340382 100872 340562 100960
rect 340670 100872 340850 100960
rect 340958 100872 341138 100960
rect 341246 100872 341426 100960
rect 341534 100872 341714 100960
rect 341822 100872 342002 100960
rect 354302 100872 354482 100960
rect 354590 100872 354770 100960
rect 354878 100872 355058 100960
rect 355166 100872 355346 100960
rect 355454 100872 355634 100960
rect 355742 100872 355922 100960
rect 356030 100872 356210 100960
rect 356318 100872 356498 100960
rect 368798 100872 368978 100960
rect 369086 100872 369266 100960
rect 369374 100872 369554 100960
rect 369662 100872 369842 100960
rect 369950 100872 370130 100960
rect 370238 100872 370418 100960
rect 370526 100872 370706 100960
rect 370814 100872 370994 100960
rect 383294 100872 383474 100960
rect 383582 100872 383762 100960
rect 383870 100872 384050 100960
rect 384158 100872 384338 100960
rect 384446 100872 384626 100960
rect 384734 100872 384914 100960
rect 385022 100872 385202 100960
rect 385310 100872 385490 100960
rect 397790 100872 397970 100960
rect 398078 100872 398258 100960
rect 398366 100872 398546 100960
rect 398654 100872 398834 100960
rect 398942 100872 399122 100960
rect 399230 100872 399410 100960
rect 399518 100872 399698 100960
rect 399806 100872 399986 100960
rect 412286 100872 412466 100960
rect 412574 100872 412754 100960
rect 412862 100872 413042 100960
rect 413150 100872 413330 100960
rect 413438 100872 413618 100960
rect 413726 100872 413906 100960
rect 414014 100872 414194 100960
rect 414302 100872 414482 100960
rect 426782 100872 426962 100960
rect 427070 100872 427250 100960
rect 427358 100872 427538 100960
rect 427646 100872 427826 100960
rect 427934 100872 428114 100960
rect 428222 100872 428402 100960
rect 428510 100872 428690 100960
rect 428798 100872 428978 100960
rect 441278 100872 441458 100960
rect 441566 100872 441746 100960
rect 441854 100872 442034 100960
rect 442142 100872 442322 100960
rect 442430 100872 442610 100960
rect 442718 100872 442898 100960
rect 443006 100872 443186 100960
rect 443294 100872 443474 100960
rect 455774 100872 455954 100960
rect 456062 100872 456242 100960
rect 456350 100872 456530 100960
rect 456638 100872 456818 100960
rect 456926 100872 457106 100960
rect 457214 100872 457394 100960
rect 457502 100872 457682 100960
rect 457790 100872 457970 100960
rect 180350 100396 180530 100484
rect 180638 100396 180818 100484
rect 180926 100396 181106 100484
rect 181214 100396 181394 100484
rect 181502 100396 181682 100484
rect 181790 100396 181970 100484
rect 182078 100396 182258 100484
rect 182366 100396 182546 100484
rect 194846 100396 195026 100484
rect 195134 100396 195314 100484
rect 195422 100396 195602 100484
rect 195710 100396 195890 100484
rect 195998 100396 196178 100484
rect 196286 100396 196466 100484
rect 196574 100396 196754 100484
rect 196862 100396 197042 100484
rect 209342 100396 209522 100484
rect 209630 100396 209810 100484
rect 209918 100396 210098 100484
rect 210206 100396 210386 100484
rect 210494 100396 210674 100484
rect 210782 100396 210962 100484
rect 211070 100396 211250 100484
rect 211358 100396 211538 100484
rect 223838 100396 224018 100484
rect 224126 100396 224306 100484
rect 224414 100396 224594 100484
rect 224702 100396 224882 100484
rect 224990 100396 225170 100484
rect 225278 100396 225458 100484
rect 225566 100396 225746 100484
rect 225854 100396 226034 100484
rect 238334 100396 238514 100484
rect 238622 100396 238802 100484
rect 238910 100396 239090 100484
rect 239198 100396 239378 100484
rect 239486 100396 239666 100484
rect 239774 100396 239954 100484
rect 240062 100396 240242 100484
rect 240350 100396 240530 100484
rect 252830 100396 253010 100484
rect 253118 100396 253298 100484
rect 253406 100396 253586 100484
rect 253694 100396 253874 100484
rect 253982 100396 254162 100484
rect 254270 100396 254450 100484
rect 254558 100396 254738 100484
rect 254846 100396 255026 100484
rect 267326 100396 267506 100484
rect 267614 100396 267794 100484
rect 267902 100396 268082 100484
rect 268190 100396 268370 100484
rect 268478 100396 268658 100484
rect 268766 100396 268946 100484
rect 269054 100396 269234 100484
rect 269342 100396 269522 100484
rect 281822 100396 282002 100484
rect 282110 100396 282290 100484
rect 282398 100396 282578 100484
rect 282686 100396 282866 100484
rect 282974 100396 283154 100484
rect 283262 100396 283442 100484
rect 283550 100396 283730 100484
rect 283838 100396 284018 100484
rect 296318 100396 296498 100484
rect 296606 100396 296786 100484
rect 296894 100396 297074 100484
rect 297182 100396 297362 100484
rect 297470 100396 297650 100484
rect 297758 100396 297938 100484
rect 298046 100396 298226 100484
rect 298334 100396 298514 100484
rect 310814 100396 310994 100484
rect 311102 100396 311282 100484
rect 311390 100396 311570 100484
rect 311678 100396 311858 100484
rect 311966 100396 312146 100484
rect 312254 100396 312434 100484
rect 312542 100396 312722 100484
rect 312830 100396 313010 100484
rect 325310 100396 325490 100484
rect 325598 100396 325778 100484
rect 325886 100396 326066 100484
rect 326174 100396 326354 100484
rect 326462 100396 326642 100484
rect 326750 100396 326930 100484
rect 327038 100396 327218 100484
rect 327326 100396 327506 100484
rect 339806 100396 339986 100484
rect 340094 100396 340274 100484
rect 340382 100396 340562 100484
rect 340670 100396 340850 100484
rect 340958 100396 341138 100484
rect 341246 100396 341426 100484
rect 341534 100396 341714 100484
rect 341822 100396 342002 100484
rect 354302 100396 354482 100484
rect 354590 100396 354770 100484
rect 354878 100396 355058 100484
rect 355166 100396 355346 100484
rect 355454 100396 355634 100484
rect 355742 100396 355922 100484
rect 356030 100396 356210 100484
rect 356318 100396 356498 100484
rect 368798 100396 368978 100484
rect 369086 100396 369266 100484
rect 369374 100396 369554 100484
rect 369662 100396 369842 100484
rect 369950 100396 370130 100484
rect 370238 100396 370418 100484
rect 370526 100396 370706 100484
rect 370814 100396 370994 100484
rect 383294 100396 383474 100484
rect 383582 100396 383762 100484
rect 383870 100396 384050 100484
rect 384158 100396 384338 100484
rect 384446 100396 384626 100484
rect 384734 100396 384914 100484
rect 385022 100396 385202 100484
rect 385310 100396 385490 100484
rect 397790 100396 397970 100484
rect 398078 100396 398258 100484
rect 398366 100396 398546 100484
rect 398654 100396 398834 100484
rect 398942 100396 399122 100484
rect 399230 100396 399410 100484
rect 399518 100396 399698 100484
rect 399806 100396 399986 100484
rect 412286 100396 412466 100484
rect 412574 100396 412754 100484
rect 412862 100396 413042 100484
rect 413150 100396 413330 100484
rect 413438 100396 413618 100484
rect 413726 100396 413906 100484
rect 414014 100396 414194 100484
rect 414302 100396 414482 100484
rect 426782 100396 426962 100484
rect 427070 100396 427250 100484
rect 427358 100396 427538 100484
rect 427646 100396 427826 100484
rect 427934 100396 428114 100484
rect 428222 100396 428402 100484
rect 428510 100396 428690 100484
rect 428798 100396 428978 100484
rect 441278 100396 441458 100484
rect 441566 100396 441746 100484
rect 441854 100396 442034 100484
rect 442142 100396 442322 100484
rect 442430 100396 442610 100484
rect 442718 100396 442898 100484
rect 443006 100396 443186 100484
rect 443294 100396 443474 100484
rect 455774 100396 455954 100484
rect 456062 100396 456242 100484
rect 456350 100396 456530 100484
rect 456638 100396 456818 100484
rect 456926 100396 457106 100484
rect 457214 100396 457394 100484
rect 457502 100396 457682 100484
rect 457790 100396 457970 100484
rect 180350 100180 180530 100268
rect 180638 100180 180818 100268
rect 180926 100180 181106 100268
rect 181214 100180 181394 100268
rect 181502 100180 181682 100268
rect 181790 100180 181970 100268
rect 182078 100180 182258 100268
rect 182366 100180 182546 100268
rect 194846 100180 195026 100268
rect 195134 100180 195314 100268
rect 195422 100180 195602 100268
rect 195710 100180 195890 100268
rect 195998 100180 196178 100268
rect 196286 100180 196466 100268
rect 196574 100180 196754 100268
rect 196862 100180 197042 100268
rect 209342 100180 209522 100268
rect 209630 100180 209810 100268
rect 209918 100180 210098 100268
rect 210206 100180 210386 100268
rect 210494 100180 210674 100268
rect 210782 100180 210962 100268
rect 211070 100180 211250 100268
rect 211358 100180 211538 100268
rect 223838 100180 224018 100268
rect 224126 100180 224306 100268
rect 224414 100180 224594 100268
rect 224702 100180 224882 100268
rect 224990 100180 225170 100268
rect 225278 100180 225458 100268
rect 225566 100180 225746 100268
rect 225854 100180 226034 100268
rect 238334 100180 238514 100268
rect 238622 100180 238802 100268
rect 238910 100180 239090 100268
rect 239198 100180 239378 100268
rect 239486 100180 239666 100268
rect 239774 100180 239954 100268
rect 240062 100180 240242 100268
rect 240350 100180 240530 100268
rect 252830 100180 253010 100268
rect 253118 100180 253298 100268
rect 253406 100180 253586 100268
rect 253694 100180 253874 100268
rect 253982 100180 254162 100268
rect 254270 100180 254450 100268
rect 254558 100180 254738 100268
rect 254846 100180 255026 100268
rect 267326 100180 267506 100268
rect 267614 100180 267794 100268
rect 267902 100180 268082 100268
rect 268190 100180 268370 100268
rect 268478 100180 268658 100268
rect 268766 100180 268946 100268
rect 269054 100180 269234 100268
rect 269342 100180 269522 100268
rect 281822 100180 282002 100268
rect 282110 100180 282290 100268
rect 282398 100180 282578 100268
rect 282686 100180 282866 100268
rect 282974 100180 283154 100268
rect 283262 100180 283442 100268
rect 283550 100180 283730 100268
rect 283838 100180 284018 100268
rect 296318 100180 296498 100268
rect 296606 100180 296786 100268
rect 296894 100180 297074 100268
rect 297182 100180 297362 100268
rect 297470 100180 297650 100268
rect 297758 100180 297938 100268
rect 298046 100180 298226 100268
rect 298334 100180 298514 100268
rect 310814 100180 310994 100268
rect 311102 100180 311282 100268
rect 311390 100180 311570 100268
rect 311678 100180 311858 100268
rect 311966 100180 312146 100268
rect 312254 100180 312434 100268
rect 312542 100180 312722 100268
rect 312830 100180 313010 100268
rect 325310 100180 325490 100268
rect 325598 100180 325778 100268
rect 325886 100180 326066 100268
rect 326174 100180 326354 100268
rect 326462 100180 326642 100268
rect 326750 100180 326930 100268
rect 327038 100180 327218 100268
rect 327326 100180 327506 100268
rect 339806 100180 339986 100268
rect 340094 100180 340274 100268
rect 340382 100180 340562 100268
rect 340670 100180 340850 100268
rect 340958 100180 341138 100268
rect 341246 100180 341426 100268
rect 341534 100180 341714 100268
rect 341822 100180 342002 100268
rect 354302 100180 354482 100268
rect 354590 100180 354770 100268
rect 354878 100180 355058 100268
rect 355166 100180 355346 100268
rect 355454 100180 355634 100268
rect 355742 100180 355922 100268
rect 356030 100180 356210 100268
rect 356318 100180 356498 100268
rect 368798 100180 368978 100268
rect 369086 100180 369266 100268
rect 369374 100180 369554 100268
rect 369662 100180 369842 100268
rect 369950 100180 370130 100268
rect 370238 100180 370418 100268
rect 370526 100180 370706 100268
rect 370814 100180 370994 100268
rect 383294 100180 383474 100268
rect 383582 100180 383762 100268
rect 383870 100180 384050 100268
rect 384158 100180 384338 100268
rect 384446 100180 384626 100268
rect 384734 100180 384914 100268
rect 385022 100180 385202 100268
rect 385310 100180 385490 100268
rect 397790 100180 397970 100268
rect 398078 100180 398258 100268
rect 398366 100180 398546 100268
rect 398654 100180 398834 100268
rect 398942 100180 399122 100268
rect 399230 100180 399410 100268
rect 399518 100180 399698 100268
rect 399806 100180 399986 100268
rect 412286 100180 412466 100268
rect 412574 100180 412754 100268
rect 412862 100180 413042 100268
rect 413150 100180 413330 100268
rect 413438 100180 413618 100268
rect 413726 100180 413906 100268
rect 414014 100180 414194 100268
rect 414302 100180 414482 100268
rect 426782 100180 426962 100268
rect 427070 100180 427250 100268
rect 427358 100180 427538 100268
rect 427646 100180 427826 100268
rect 427934 100180 428114 100268
rect 428222 100180 428402 100268
rect 428510 100180 428690 100268
rect 428798 100180 428978 100268
rect 441278 100180 441458 100268
rect 441566 100180 441746 100268
rect 441854 100180 442034 100268
rect 442142 100180 442322 100268
rect 442430 100180 442610 100268
rect 442718 100180 442898 100268
rect 443006 100180 443186 100268
rect 443294 100180 443474 100268
rect 455774 100180 455954 100268
rect 456062 100180 456242 100268
rect 456350 100180 456530 100268
rect 456638 100180 456818 100268
rect 456926 100180 457106 100268
rect 457214 100180 457394 100268
rect 457502 100180 457682 100268
rect 457790 100180 457970 100268
rect 180350 86028 180530 86116
rect 180638 86028 180818 86116
rect 180926 86028 181106 86116
rect 181214 86028 181394 86116
rect 181502 86028 181682 86116
rect 181790 86028 181970 86116
rect 182078 86028 182258 86116
rect 182366 86028 182546 86116
rect 194846 86028 195026 86116
rect 195134 86028 195314 86116
rect 195422 86028 195602 86116
rect 195710 86028 195890 86116
rect 195998 86028 196178 86116
rect 196286 86028 196466 86116
rect 196574 86028 196754 86116
rect 196862 86028 197042 86116
rect 209342 86028 209522 86116
rect 209630 86028 209810 86116
rect 209918 86028 210098 86116
rect 210206 86028 210386 86116
rect 210494 86028 210674 86116
rect 210782 86028 210962 86116
rect 211070 86028 211250 86116
rect 211358 86028 211538 86116
rect 223838 86028 224018 86116
rect 224126 86028 224306 86116
rect 224414 86028 224594 86116
rect 224702 86028 224882 86116
rect 224990 86028 225170 86116
rect 225278 86028 225458 86116
rect 225566 86028 225746 86116
rect 225854 86028 226034 86116
rect 238334 86028 238514 86116
rect 238622 86028 238802 86116
rect 238910 86028 239090 86116
rect 239198 86028 239378 86116
rect 239486 86028 239666 86116
rect 239774 86028 239954 86116
rect 240062 86028 240242 86116
rect 240350 86028 240530 86116
rect 252830 86028 253010 86116
rect 253118 86028 253298 86116
rect 253406 86028 253586 86116
rect 253694 86028 253874 86116
rect 253982 86028 254162 86116
rect 254270 86028 254450 86116
rect 254558 86028 254738 86116
rect 254846 86028 255026 86116
rect 267326 86028 267506 86116
rect 267614 86028 267794 86116
rect 267902 86028 268082 86116
rect 268190 86028 268370 86116
rect 268478 86028 268658 86116
rect 268766 86028 268946 86116
rect 269054 86028 269234 86116
rect 269342 86028 269522 86116
rect 281822 86028 282002 86116
rect 282110 86028 282290 86116
rect 282398 86028 282578 86116
rect 282686 86028 282866 86116
rect 282974 86028 283154 86116
rect 283262 86028 283442 86116
rect 283550 86028 283730 86116
rect 283838 86028 284018 86116
rect 296318 86028 296498 86116
rect 296606 86028 296786 86116
rect 296894 86028 297074 86116
rect 297182 86028 297362 86116
rect 297470 86028 297650 86116
rect 297758 86028 297938 86116
rect 298046 86028 298226 86116
rect 298334 86028 298514 86116
rect 310814 86028 310994 86116
rect 311102 86028 311282 86116
rect 311390 86028 311570 86116
rect 311678 86028 311858 86116
rect 311966 86028 312146 86116
rect 312254 86028 312434 86116
rect 312542 86028 312722 86116
rect 312830 86028 313010 86116
rect 325310 86028 325490 86116
rect 325598 86028 325778 86116
rect 325886 86028 326066 86116
rect 326174 86028 326354 86116
rect 326462 86028 326642 86116
rect 326750 86028 326930 86116
rect 327038 86028 327218 86116
rect 327326 86028 327506 86116
rect 339806 86028 339986 86116
rect 340094 86028 340274 86116
rect 340382 86028 340562 86116
rect 340670 86028 340850 86116
rect 340958 86028 341138 86116
rect 341246 86028 341426 86116
rect 341534 86028 341714 86116
rect 341822 86028 342002 86116
rect 354302 86028 354482 86116
rect 354590 86028 354770 86116
rect 354878 86028 355058 86116
rect 355166 86028 355346 86116
rect 355454 86028 355634 86116
rect 355742 86028 355922 86116
rect 356030 86028 356210 86116
rect 356318 86028 356498 86116
rect 368798 86028 368978 86116
rect 369086 86028 369266 86116
rect 369374 86028 369554 86116
rect 369662 86028 369842 86116
rect 369950 86028 370130 86116
rect 370238 86028 370418 86116
rect 370526 86028 370706 86116
rect 370814 86028 370994 86116
rect 383294 86028 383474 86116
rect 383582 86028 383762 86116
rect 383870 86028 384050 86116
rect 384158 86028 384338 86116
rect 384446 86028 384626 86116
rect 384734 86028 384914 86116
rect 385022 86028 385202 86116
rect 385310 86028 385490 86116
rect 397790 86028 397970 86116
rect 398078 86028 398258 86116
rect 398366 86028 398546 86116
rect 398654 86028 398834 86116
rect 398942 86028 399122 86116
rect 399230 86028 399410 86116
rect 399518 86028 399698 86116
rect 399806 86028 399986 86116
rect 412286 86028 412466 86116
rect 412574 86028 412754 86116
rect 412862 86028 413042 86116
rect 413150 86028 413330 86116
rect 413438 86028 413618 86116
rect 413726 86028 413906 86116
rect 414014 86028 414194 86116
rect 414302 86028 414482 86116
rect 426782 86028 426962 86116
rect 427070 86028 427250 86116
rect 427358 86028 427538 86116
rect 427646 86028 427826 86116
rect 427934 86028 428114 86116
rect 428222 86028 428402 86116
rect 428510 86028 428690 86116
rect 428798 86028 428978 86116
rect 441278 86028 441458 86116
rect 441566 86028 441746 86116
rect 441854 86028 442034 86116
rect 442142 86028 442322 86116
rect 442430 86028 442610 86116
rect 442718 86028 442898 86116
rect 443006 86028 443186 86116
rect 443294 86028 443474 86116
rect 455774 86028 455954 86116
rect 456062 86028 456242 86116
rect 456350 86028 456530 86116
rect 456638 86028 456818 86116
rect 456926 86028 457106 86116
rect 457214 86028 457394 86116
rect 457502 86028 457682 86116
rect 457790 86028 457970 86116
rect 180350 85812 180530 85900
rect 180638 85812 180818 85900
rect 180926 85812 181106 85900
rect 181214 85812 181394 85900
rect 181502 85812 181682 85900
rect 181790 85812 181970 85900
rect 182078 85812 182258 85900
rect 182366 85812 182546 85900
rect 194846 85812 195026 85900
rect 195134 85812 195314 85900
rect 195422 85812 195602 85900
rect 195710 85812 195890 85900
rect 195998 85812 196178 85900
rect 196286 85812 196466 85900
rect 196574 85812 196754 85900
rect 196862 85812 197042 85900
rect 209342 85812 209522 85900
rect 209630 85812 209810 85900
rect 209918 85812 210098 85900
rect 210206 85812 210386 85900
rect 210494 85812 210674 85900
rect 210782 85812 210962 85900
rect 211070 85812 211250 85900
rect 211358 85812 211538 85900
rect 223838 85812 224018 85900
rect 224126 85812 224306 85900
rect 224414 85812 224594 85900
rect 224702 85812 224882 85900
rect 224990 85812 225170 85900
rect 225278 85812 225458 85900
rect 225566 85812 225746 85900
rect 225854 85812 226034 85900
rect 238334 85812 238514 85900
rect 238622 85812 238802 85900
rect 238910 85812 239090 85900
rect 239198 85812 239378 85900
rect 239486 85812 239666 85900
rect 239774 85812 239954 85900
rect 240062 85812 240242 85900
rect 240350 85812 240530 85900
rect 252830 85812 253010 85900
rect 253118 85812 253298 85900
rect 253406 85812 253586 85900
rect 253694 85812 253874 85900
rect 253982 85812 254162 85900
rect 254270 85812 254450 85900
rect 254558 85812 254738 85900
rect 254846 85812 255026 85900
rect 267326 85812 267506 85900
rect 267614 85812 267794 85900
rect 267902 85812 268082 85900
rect 268190 85812 268370 85900
rect 268478 85812 268658 85900
rect 268766 85812 268946 85900
rect 269054 85812 269234 85900
rect 269342 85812 269522 85900
rect 281822 85812 282002 85900
rect 282110 85812 282290 85900
rect 282398 85812 282578 85900
rect 282686 85812 282866 85900
rect 282974 85812 283154 85900
rect 283262 85812 283442 85900
rect 283550 85812 283730 85900
rect 283838 85812 284018 85900
rect 296318 85812 296498 85900
rect 296606 85812 296786 85900
rect 296894 85812 297074 85900
rect 297182 85812 297362 85900
rect 297470 85812 297650 85900
rect 297758 85812 297938 85900
rect 298046 85812 298226 85900
rect 298334 85812 298514 85900
rect 310814 85812 310994 85900
rect 311102 85812 311282 85900
rect 311390 85812 311570 85900
rect 311678 85812 311858 85900
rect 311966 85812 312146 85900
rect 312254 85812 312434 85900
rect 312542 85812 312722 85900
rect 312830 85812 313010 85900
rect 325310 85812 325490 85900
rect 325598 85812 325778 85900
rect 325886 85812 326066 85900
rect 326174 85812 326354 85900
rect 326462 85812 326642 85900
rect 326750 85812 326930 85900
rect 327038 85812 327218 85900
rect 327326 85812 327506 85900
rect 339806 85812 339986 85900
rect 340094 85812 340274 85900
rect 340382 85812 340562 85900
rect 340670 85812 340850 85900
rect 340958 85812 341138 85900
rect 341246 85812 341426 85900
rect 341534 85812 341714 85900
rect 341822 85812 342002 85900
rect 354302 85812 354482 85900
rect 354590 85812 354770 85900
rect 354878 85812 355058 85900
rect 355166 85812 355346 85900
rect 355454 85812 355634 85900
rect 355742 85812 355922 85900
rect 356030 85812 356210 85900
rect 356318 85812 356498 85900
rect 368798 85812 368978 85900
rect 369086 85812 369266 85900
rect 369374 85812 369554 85900
rect 369662 85812 369842 85900
rect 369950 85812 370130 85900
rect 370238 85812 370418 85900
rect 370526 85812 370706 85900
rect 370814 85812 370994 85900
rect 383294 85812 383474 85900
rect 383582 85812 383762 85900
rect 383870 85812 384050 85900
rect 384158 85812 384338 85900
rect 384446 85812 384626 85900
rect 384734 85812 384914 85900
rect 385022 85812 385202 85900
rect 385310 85812 385490 85900
rect 397790 85812 397970 85900
rect 398078 85812 398258 85900
rect 398366 85812 398546 85900
rect 398654 85812 398834 85900
rect 398942 85812 399122 85900
rect 399230 85812 399410 85900
rect 399518 85812 399698 85900
rect 399806 85812 399986 85900
rect 412286 85812 412466 85900
rect 412574 85812 412754 85900
rect 412862 85812 413042 85900
rect 413150 85812 413330 85900
rect 413438 85812 413618 85900
rect 413726 85812 413906 85900
rect 414014 85812 414194 85900
rect 414302 85812 414482 85900
rect 426782 85812 426962 85900
rect 427070 85812 427250 85900
rect 427358 85812 427538 85900
rect 427646 85812 427826 85900
rect 427934 85812 428114 85900
rect 428222 85812 428402 85900
rect 428510 85812 428690 85900
rect 428798 85812 428978 85900
rect 441278 85812 441458 85900
rect 441566 85812 441746 85900
rect 441854 85812 442034 85900
rect 442142 85812 442322 85900
rect 442430 85812 442610 85900
rect 442718 85812 442898 85900
rect 443006 85812 443186 85900
rect 443294 85812 443474 85900
rect 455774 85812 455954 85900
rect 456062 85812 456242 85900
rect 456350 85812 456530 85900
rect 456638 85812 456818 85900
rect 456926 85812 457106 85900
rect 457214 85812 457394 85900
rect 457502 85812 457682 85900
rect 457790 85812 457970 85900
rect 180350 85336 180530 85424
rect 180638 85336 180818 85424
rect 180926 85336 181106 85424
rect 181214 85336 181394 85424
rect 181502 85336 181682 85424
rect 181790 85336 181970 85424
rect 182078 85336 182258 85424
rect 182366 85336 182546 85424
rect 194846 85336 195026 85424
rect 195134 85336 195314 85424
rect 195422 85336 195602 85424
rect 195710 85336 195890 85424
rect 195998 85336 196178 85424
rect 196286 85336 196466 85424
rect 196574 85336 196754 85424
rect 196862 85336 197042 85424
rect 209342 85336 209522 85424
rect 209630 85336 209810 85424
rect 209918 85336 210098 85424
rect 210206 85336 210386 85424
rect 210494 85336 210674 85424
rect 210782 85336 210962 85424
rect 211070 85336 211250 85424
rect 211358 85336 211538 85424
rect 223838 85336 224018 85424
rect 224126 85336 224306 85424
rect 224414 85336 224594 85424
rect 224702 85336 224882 85424
rect 224990 85336 225170 85424
rect 225278 85336 225458 85424
rect 225566 85336 225746 85424
rect 225854 85336 226034 85424
rect 238334 85336 238514 85424
rect 238622 85336 238802 85424
rect 238910 85336 239090 85424
rect 239198 85336 239378 85424
rect 239486 85336 239666 85424
rect 239774 85336 239954 85424
rect 240062 85336 240242 85424
rect 240350 85336 240530 85424
rect 252830 85336 253010 85424
rect 253118 85336 253298 85424
rect 253406 85336 253586 85424
rect 253694 85336 253874 85424
rect 253982 85336 254162 85424
rect 254270 85336 254450 85424
rect 254558 85336 254738 85424
rect 254846 85336 255026 85424
rect 267326 85336 267506 85424
rect 267614 85336 267794 85424
rect 267902 85336 268082 85424
rect 268190 85336 268370 85424
rect 268478 85336 268658 85424
rect 268766 85336 268946 85424
rect 269054 85336 269234 85424
rect 269342 85336 269522 85424
rect 281822 85336 282002 85424
rect 282110 85336 282290 85424
rect 282398 85336 282578 85424
rect 282686 85336 282866 85424
rect 282974 85336 283154 85424
rect 283262 85336 283442 85424
rect 283550 85336 283730 85424
rect 283838 85336 284018 85424
rect 296318 85336 296498 85424
rect 296606 85336 296786 85424
rect 296894 85336 297074 85424
rect 297182 85336 297362 85424
rect 297470 85336 297650 85424
rect 297758 85336 297938 85424
rect 298046 85336 298226 85424
rect 298334 85336 298514 85424
rect 310814 85336 310994 85424
rect 311102 85336 311282 85424
rect 311390 85336 311570 85424
rect 311678 85336 311858 85424
rect 311966 85336 312146 85424
rect 312254 85336 312434 85424
rect 312542 85336 312722 85424
rect 312830 85336 313010 85424
rect 325310 85336 325490 85424
rect 325598 85336 325778 85424
rect 325886 85336 326066 85424
rect 326174 85336 326354 85424
rect 326462 85336 326642 85424
rect 326750 85336 326930 85424
rect 327038 85336 327218 85424
rect 327326 85336 327506 85424
rect 339806 85336 339986 85424
rect 340094 85336 340274 85424
rect 340382 85336 340562 85424
rect 340670 85336 340850 85424
rect 340958 85336 341138 85424
rect 341246 85336 341426 85424
rect 341534 85336 341714 85424
rect 341822 85336 342002 85424
rect 354302 85336 354482 85424
rect 354590 85336 354770 85424
rect 354878 85336 355058 85424
rect 355166 85336 355346 85424
rect 355454 85336 355634 85424
rect 355742 85336 355922 85424
rect 356030 85336 356210 85424
rect 356318 85336 356498 85424
rect 368798 85336 368978 85424
rect 369086 85336 369266 85424
rect 369374 85336 369554 85424
rect 369662 85336 369842 85424
rect 369950 85336 370130 85424
rect 370238 85336 370418 85424
rect 370526 85336 370706 85424
rect 370814 85336 370994 85424
rect 383294 85336 383474 85424
rect 383582 85336 383762 85424
rect 383870 85336 384050 85424
rect 384158 85336 384338 85424
rect 384446 85336 384626 85424
rect 384734 85336 384914 85424
rect 385022 85336 385202 85424
rect 385310 85336 385490 85424
rect 397790 85336 397970 85424
rect 398078 85336 398258 85424
rect 398366 85336 398546 85424
rect 398654 85336 398834 85424
rect 398942 85336 399122 85424
rect 399230 85336 399410 85424
rect 399518 85336 399698 85424
rect 399806 85336 399986 85424
rect 412286 85336 412466 85424
rect 412574 85336 412754 85424
rect 412862 85336 413042 85424
rect 413150 85336 413330 85424
rect 413438 85336 413618 85424
rect 413726 85336 413906 85424
rect 414014 85336 414194 85424
rect 414302 85336 414482 85424
rect 426782 85336 426962 85424
rect 427070 85336 427250 85424
rect 427358 85336 427538 85424
rect 427646 85336 427826 85424
rect 427934 85336 428114 85424
rect 428222 85336 428402 85424
rect 428510 85336 428690 85424
rect 428798 85336 428978 85424
rect 441278 85336 441458 85424
rect 441566 85336 441746 85424
rect 441854 85336 442034 85424
rect 442142 85336 442322 85424
rect 442430 85336 442610 85424
rect 442718 85336 442898 85424
rect 443006 85336 443186 85424
rect 443294 85336 443474 85424
rect 455774 85336 455954 85424
rect 456062 85336 456242 85424
rect 456350 85336 456530 85424
rect 456638 85336 456818 85424
rect 456926 85336 457106 85424
rect 457214 85336 457394 85424
rect 457502 85336 457682 85424
rect 457790 85336 457970 85424
rect 180350 85120 180530 85208
rect 180638 85120 180818 85208
rect 180926 85120 181106 85208
rect 181214 85120 181394 85208
rect 181502 85120 181682 85208
rect 181790 85120 181970 85208
rect 182078 85120 182258 85208
rect 182366 85120 182546 85208
rect 194846 85120 195026 85208
rect 195134 85120 195314 85208
rect 195422 85120 195602 85208
rect 195710 85120 195890 85208
rect 195998 85120 196178 85208
rect 196286 85120 196466 85208
rect 196574 85120 196754 85208
rect 196862 85120 197042 85208
rect 209342 85120 209522 85208
rect 209630 85120 209810 85208
rect 209918 85120 210098 85208
rect 210206 85120 210386 85208
rect 210494 85120 210674 85208
rect 210782 85120 210962 85208
rect 211070 85120 211250 85208
rect 211358 85120 211538 85208
rect 223838 85120 224018 85208
rect 224126 85120 224306 85208
rect 224414 85120 224594 85208
rect 224702 85120 224882 85208
rect 224990 85120 225170 85208
rect 225278 85120 225458 85208
rect 225566 85120 225746 85208
rect 225854 85120 226034 85208
rect 238334 85120 238514 85208
rect 238622 85120 238802 85208
rect 238910 85120 239090 85208
rect 239198 85120 239378 85208
rect 239486 85120 239666 85208
rect 239774 85120 239954 85208
rect 240062 85120 240242 85208
rect 240350 85120 240530 85208
rect 252830 85120 253010 85208
rect 253118 85120 253298 85208
rect 253406 85120 253586 85208
rect 253694 85120 253874 85208
rect 253982 85120 254162 85208
rect 254270 85120 254450 85208
rect 254558 85120 254738 85208
rect 254846 85120 255026 85208
rect 267326 85120 267506 85208
rect 267614 85120 267794 85208
rect 267902 85120 268082 85208
rect 268190 85120 268370 85208
rect 268478 85120 268658 85208
rect 268766 85120 268946 85208
rect 269054 85120 269234 85208
rect 269342 85120 269522 85208
rect 281822 85120 282002 85208
rect 282110 85120 282290 85208
rect 282398 85120 282578 85208
rect 282686 85120 282866 85208
rect 282974 85120 283154 85208
rect 283262 85120 283442 85208
rect 283550 85120 283730 85208
rect 283838 85120 284018 85208
rect 296318 85120 296498 85208
rect 296606 85120 296786 85208
rect 296894 85120 297074 85208
rect 297182 85120 297362 85208
rect 297470 85120 297650 85208
rect 297758 85120 297938 85208
rect 298046 85120 298226 85208
rect 298334 85120 298514 85208
rect 310814 85120 310994 85208
rect 311102 85120 311282 85208
rect 311390 85120 311570 85208
rect 311678 85120 311858 85208
rect 311966 85120 312146 85208
rect 312254 85120 312434 85208
rect 312542 85120 312722 85208
rect 312830 85120 313010 85208
rect 325310 85120 325490 85208
rect 325598 85120 325778 85208
rect 325886 85120 326066 85208
rect 326174 85120 326354 85208
rect 326462 85120 326642 85208
rect 326750 85120 326930 85208
rect 327038 85120 327218 85208
rect 327326 85120 327506 85208
rect 339806 85120 339986 85208
rect 340094 85120 340274 85208
rect 340382 85120 340562 85208
rect 340670 85120 340850 85208
rect 340958 85120 341138 85208
rect 341246 85120 341426 85208
rect 341534 85120 341714 85208
rect 341822 85120 342002 85208
rect 354302 85120 354482 85208
rect 354590 85120 354770 85208
rect 354878 85120 355058 85208
rect 355166 85120 355346 85208
rect 355454 85120 355634 85208
rect 355742 85120 355922 85208
rect 356030 85120 356210 85208
rect 356318 85120 356498 85208
rect 368798 85120 368978 85208
rect 369086 85120 369266 85208
rect 369374 85120 369554 85208
rect 369662 85120 369842 85208
rect 369950 85120 370130 85208
rect 370238 85120 370418 85208
rect 370526 85120 370706 85208
rect 370814 85120 370994 85208
rect 383294 85120 383474 85208
rect 383582 85120 383762 85208
rect 383870 85120 384050 85208
rect 384158 85120 384338 85208
rect 384446 85120 384626 85208
rect 384734 85120 384914 85208
rect 385022 85120 385202 85208
rect 385310 85120 385490 85208
rect 397790 85120 397970 85208
rect 398078 85120 398258 85208
rect 398366 85120 398546 85208
rect 398654 85120 398834 85208
rect 398942 85120 399122 85208
rect 399230 85120 399410 85208
rect 399518 85120 399698 85208
rect 399806 85120 399986 85208
rect 412286 85120 412466 85208
rect 412574 85120 412754 85208
rect 412862 85120 413042 85208
rect 413150 85120 413330 85208
rect 413438 85120 413618 85208
rect 413726 85120 413906 85208
rect 414014 85120 414194 85208
rect 414302 85120 414482 85208
rect 426782 85120 426962 85208
rect 427070 85120 427250 85208
rect 427358 85120 427538 85208
rect 427646 85120 427826 85208
rect 427934 85120 428114 85208
rect 428222 85120 428402 85208
rect 428510 85120 428690 85208
rect 428798 85120 428978 85208
rect 441278 85120 441458 85208
rect 441566 85120 441746 85208
rect 441854 85120 442034 85208
rect 442142 85120 442322 85208
rect 442430 85120 442610 85208
rect 442718 85120 442898 85208
rect 443006 85120 443186 85208
rect 443294 85120 443474 85208
rect 455774 85120 455954 85208
rect 456062 85120 456242 85208
rect 456350 85120 456530 85208
rect 456638 85120 456818 85208
rect 456926 85120 457106 85208
rect 457214 85120 457394 85208
rect 457502 85120 457682 85208
rect 457790 85120 457970 85208
rect 180350 70968 180530 71056
rect 180638 70968 180818 71056
rect 180926 70968 181106 71056
rect 181214 70968 181394 71056
rect 181502 70968 181682 71056
rect 181790 70968 181970 71056
rect 182078 70968 182258 71056
rect 182366 70968 182546 71056
rect 194846 70968 195026 71056
rect 195134 70968 195314 71056
rect 195422 70968 195602 71056
rect 195710 70968 195890 71056
rect 195998 70968 196178 71056
rect 196286 70968 196466 71056
rect 196574 70968 196754 71056
rect 196862 70968 197042 71056
rect 209342 70968 209522 71056
rect 209630 70968 209810 71056
rect 209918 70968 210098 71056
rect 210206 70968 210386 71056
rect 210494 70968 210674 71056
rect 210782 70968 210962 71056
rect 211070 70968 211250 71056
rect 211358 70968 211538 71056
rect 223838 70968 224018 71056
rect 224126 70968 224306 71056
rect 224414 70968 224594 71056
rect 224702 70968 224882 71056
rect 224990 70968 225170 71056
rect 225278 70968 225458 71056
rect 225566 70968 225746 71056
rect 225854 70968 226034 71056
rect 238334 70968 238514 71056
rect 238622 70968 238802 71056
rect 238910 70968 239090 71056
rect 239198 70968 239378 71056
rect 239486 70968 239666 71056
rect 239774 70968 239954 71056
rect 240062 70968 240242 71056
rect 240350 70968 240530 71056
rect 252830 70968 253010 71056
rect 253118 70968 253298 71056
rect 253406 70968 253586 71056
rect 253694 70968 253874 71056
rect 253982 70968 254162 71056
rect 254270 70968 254450 71056
rect 254558 70968 254738 71056
rect 254846 70968 255026 71056
rect 267326 70968 267506 71056
rect 267614 70968 267794 71056
rect 267902 70968 268082 71056
rect 268190 70968 268370 71056
rect 268478 70968 268658 71056
rect 268766 70968 268946 71056
rect 269054 70968 269234 71056
rect 269342 70968 269522 71056
rect 281822 70968 282002 71056
rect 282110 70968 282290 71056
rect 282398 70968 282578 71056
rect 282686 70968 282866 71056
rect 282974 70968 283154 71056
rect 283262 70968 283442 71056
rect 283550 70968 283730 71056
rect 283838 70968 284018 71056
rect 296318 70968 296498 71056
rect 296606 70968 296786 71056
rect 296894 70968 297074 71056
rect 297182 70968 297362 71056
rect 297470 70968 297650 71056
rect 297758 70968 297938 71056
rect 298046 70968 298226 71056
rect 298334 70968 298514 71056
rect 310814 70968 310994 71056
rect 311102 70968 311282 71056
rect 311390 70968 311570 71056
rect 311678 70968 311858 71056
rect 311966 70968 312146 71056
rect 312254 70968 312434 71056
rect 312542 70968 312722 71056
rect 312830 70968 313010 71056
rect 325310 70968 325490 71056
rect 325598 70968 325778 71056
rect 325886 70968 326066 71056
rect 326174 70968 326354 71056
rect 326462 70968 326642 71056
rect 326750 70968 326930 71056
rect 327038 70968 327218 71056
rect 327326 70968 327506 71056
rect 339806 70968 339986 71056
rect 340094 70968 340274 71056
rect 340382 70968 340562 71056
rect 340670 70968 340850 71056
rect 340958 70968 341138 71056
rect 341246 70968 341426 71056
rect 341534 70968 341714 71056
rect 341822 70968 342002 71056
rect 354302 70968 354482 71056
rect 354590 70968 354770 71056
rect 354878 70968 355058 71056
rect 355166 70968 355346 71056
rect 355454 70968 355634 71056
rect 355742 70968 355922 71056
rect 356030 70968 356210 71056
rect 356318 70968 356498 71056
rect 368798 70968 368978 71056
rect 369086 70968 369266 71056
rect 369374 70968 369554 71056
rect 369662 70968 369842 71056
rect 369950 70968 370130 71056
rect 370238 70968 370418 71056
rect 370526 70968 370706 71056
rect 370814 70968 370994 71056
rect 383294 70968 383474 71056
rect 383582 70968 383762 71056
rect 383870 70968 384050 71056
rect 384158 70968 384338 71056
rect 384446 70968 384626 71056
rect 384734 70968 384914 71056
rect 385022 70968 385202 71056
rect 385310 70968 385490 71056
rect 397790 70968 397970 71056
rect 398078 70968 398258 71056
rect 398366 70968 398546 71056
rect 398654 70968 398834 71056
rect 398942 70968 399122 71056
rect 399230 70968 399410 71056
rect 399518 70968 399698 71056
rect 399806 70968 399986 71056
rect 412286 70968 412466 71056
rect 412574 70968 412754 71056
rect 412862 70968 413042 71056
rect 413150 70968 413330 71056
rect 413438 70968 413618 71056
rect 413726 70968 413906 71056
rect 414014 70968 414194 71056
rect 414302 70968 414482 71056
rect 426782 70968 426962 71056
rect 427070 70968 427250 71056
rect 427358 70968 427538 71056
rect 427646 70968 427826 71056
rect 427934 70968 428114 71056
rect 428222 70968 428402 71056
rect 428510 70968 428690 71056
rect 428798 70968 428978 71056
rect 441278 70968 441458 71056
rect 441566 70968 441746 71056
rect 441854 70968 442034 71056
rect 442142 70968 442322 71056
rect 442430 70968 442610 71056
rect 442718 70968 442898 71056
rect 443006 70968 443186 71056
rect 443294 70968 443474 71056
rect 455774 70968 455954 71056
rect 456062 70968 456242 71056
rect 456350 70968 456530 71056
rect 456638 70968 456818 71056
rect 456926 70968 457106 71056
rect 457214 70968 457394 71056
rect 457502 70968 457682 71056
rect 457790 70968 457970 71056
rect 180350 70752 180530 70840
rect 180638 70752 180818 70840
rect 180926 70752 181106 70840
rect 181214 70752 181394 70840
rect 181502 70752 181682 70840
rect 181790 70752 181970 70840
rect 182078 70752 182258 70840
rect 182366 70752 182546 70840
rect 194846 70752 195026 70840
rect 195134 70752 195314 70840
rect 195422 70752 195602 70840
rect 195710 70752 195890 70840
rect 195998 70752 196178 70840
rect 196286 70752 196466 70840
rect 196574 70752 196754 70840
rect 196862 70752 197042 70840
rect 209342 70752 209522 70840
rect 209630 70752 209810 70840
rect 209918 70752 210098 70840
rect 210206 70752 210386 70840
rect 210494 70752 210674 70840
rect 210782 70752 210962 70840
rect 211070 70752 211250 70840
rect 211358 70752 211538 70840
rect 223838 70752 224018 70840
rect 224126 70752 224306 70840
rect 224414 70752 224594 70840
rect 224702 70752 224882 70840
rect 224990 70752 225170 70840
rect 225278 70752 225458 70840
rect 225566 70752 225746 70840
rect 225854 70752 226034 70840
rect 238334 70752 238514 70840
rect 238622 70752 238802 70840
rect 238910 70752 239090 70840
rect 239198 70752 239378 70840
rect 239486 70752 239666 70840
rect 239774 70752 239954 70840
rect 240062 70752 240242 70840
rect 240350 70752 240530 70840
rect 252830 70752 253010 70840
rect 253118 70752 253298 70840
rect 253406 70752 253586 70840
rect 253694 70752 253874 70840
rect 253982 70752 254162 70840
rect 254270 70752 254450 70840
rect 254558 70752 254738 70840
rect 254846 70752 255026 70840
rect 267326 70752 267506 70840
rect 267614 70752 267794 70840
rect 267902 70752 268082 70840
rect 268190 70752 268370 70840
rect 268478 70752 268658 70840
rect 268766 70752 268946 70840
rect 269054 70752 269234 70840
rect 269342 70752 269522 70840
rect 281822 70752 282002 70840
rect 282110 70752 282290 70840
rect 282398 70752 282578 70840
rect 282686 70752 282866 70840
rect 282974 70752 283154 70840
rect 283262 70752 283442 70840
rect 283550 70752 283730 70840
rect 283838 70752 284018 70840
rect 296318 70752 296498 70840
rect 296606 70752 296786 70840
rect 296894 70752 297074 70840
rect 297182 70752 297362 70840
rect 297470 70752 297650 70840
rect 297758 70752 297938 70840
rect 298046 70752 298226 70840
rect 298334 70752 298514 70840
rect 310814 70752 310994 70840
rect 311102 70752 311282 70840
rect 311390 70752 311570 70840
rect 311678 70752 311858 70840
rect 311966 70752 312146 70840
rect 312254 70752 312434 70840
rect 312542 70752 312722 70840
rect 312830 70752 313010 70840
rect 325310 70752 325490 70840
rect 325598 70752 325778 70840
rect 325886 70752 326066 70840
rect 326174 70752 326354 70840
rect 326462 70752 326642 70840
rect 326750 70752 326930 70840
rect 327038 70752 327218 70840
rect 327326 70752 327506 70840
rect 339806 70752 339986 70840
rect 340094 70752 340274 70840
rect 340382 70752 340562 70840
rect 340670 70752 340850 70840
rect 340958 70752 341138 70840
rect 341246 70752 341426 70840
rect 341534 70752 341714 70840
rect 341822 70752 342002 70840
rect 354302 70752 354482 70840
rect 354590 70752 354770 70840
rect 354878 70752 355058 70840
rect 355166 70752 355346 70840
rect 355454 70752 355634 70840
rect 355742 70752 355922 70840
rect 356030 70752 356210 70840
rect 356318 70752 356498 70840
rect 368798 70752 368978 70840
rect 369086 70752 369266 70840
rect 369374 70752 369554 70840
rect 369662 70752 369842 70840
rect 369950 70752 370130 70840
rect 370238 70752 370418 70840
rect 370526 70752 370706 70840
rect 370814 70752 370994 70840
rect 383294 70752 383474 70840
rect 383582 70752 383762 70840
rect 383870 70752 384050 70840
rect 384158 70752 384338 70840
rect 384446 70752 384626 70840
rect 384734 70752 384914 70840
rect 385022 70752 385202 70840
rect 385310 70752 385490 70840
rect 397790 70752 397970 70840
rect 398078 70752 398258 70840
rect 398366 70752 398546 70840
rect 398654 70752 398834 70840
rect 398942 70752 399122 70840
rect 399230 70752 399410 70840
rect 399518 70752 399698 70840
rect 399806 70752 399986 70840
rect 412286 70752 412466 70840
rect 412574 70752 412754 70840
rect 412862 70752 413042 70840
rect 413150 70752 413330 70840
rect 413438 70752 413618 70840
rect 413726 70752 413906 70840
rect 414014 70752 414194 70840
rect 414302 70752 414482 70840
rect 426782 70752 426962 70840
rect 427070 70752 427250 70840
rect 427358 70752 427538 70840
rect 427646 70752 427826 70840
rect 427934 70752 428114 70840
rect 428222 70752 428402 70840
rect 428510 70752 428690 70840
rect 428798 70752 428978 70840
rect 441278 70752 441458 70840
rect 441566 70752 441746 70840
rect 441854 70752 442034 70840
rect 442142 70752 442322 70840
rect 442430 70752 442610 70840
rect 442718 70752 442898 70840
rect 443006 70752 443186 70840
rect 443294 70752 443474 70840
rect 455774 70752 455954 70840
rect 456062 70752 456242 70840
rect 456350 70752 456530 70840
rect 456638 70752 456818 70840
rect 456926 70752 457106 70840
rect 457214 70752 457394 70840
rect 457502 70752 457682 70840
rect 457790 70752 457970 70840
rect 180350 70276 180530 70364
rect 180638 70276 180818 70364
rect 180926 70276 181106 70364
rect 181214 70276 181394 70364
rect 181502 70276 181682 70364
rect 181790 70276 181970 70364
rect 182078 70276 182258 70364
rect 182366 70276 182546 70364
rect 194846 70276 195026 70364
rect 195134 70276 195314 70364
rect 195422 70276 195602 70364
rect 195710 70276 195890 70364
rect 195998 70276 196178 70364
rect 196286 70276 196466 70364
rect 196574 70276 196754 70364
rect 196862 70276 197042 70364
rect 209342 70276 209522 70364
rect 209630 70276 209810 70364
rect 209918 70276 210098 70364
rect 210206 70276 210386 70364
rect 210494 70276 210674 70364
rect 210782 70276 210962 70364
rect 211070 70276 211250 70364
rect 211358 70276 211538 70364
rect 223838 70276 224018 70364
rect 224126 70276 224306 70364
rect 224414 70276 224594 70364
rect 224702 70276 224882 70364
rect 224990 70276 225170 70364
rect 225278 70276 225458 70364
rect 225566 70276 225746 70364
rect 225854 70276 226034 70364
rect 238334 70276 238514 70364
rect 238622 70276 238802 70364
rect 238910 70276 239090 70364
rect 239198 70276 239378 70364
rect 239486 70276 239666 70364
rect 239774 70276 239954 70364
rect 240062 70276 240242 70364
rect 240350 70276 240530 70364
rect 252830 70276 253010 70364
rect 253118 70276 253298 70364
rect 253406 70276 253586 70364
rect 253694 70276 253874 70364
rect 253982 70276 254162 70364
rect 254270 70276 254450 70364
rect 254558 70276 254738 70364
rect 254846 70276 255026 70364
rect 267326 70276 267506 70364
rect 267614 70276 267794 70364
rect 267902 70276 268082 70364
rect 268190 70276 268370 70364
rect 268478 70276 268658 70364
rect 268766 70276 268946 70364
rect 269054 70276 269234 70364
rect 269342 70276 269522 70364
rect 281822 70276 282002 70364
rect 282110 70276 282290 70364
rect 282398 70276 282578 70364
rect 282686 70276 282866 70364
rect 282974 70276 283154 70364
rect 283262 70276 283442 70364
rect 283550 70276 283730 70364
rect 283838 70276 284018 70364
rect 296318 70276 296498 70364
rect 296606 70276 296786 70364
rect 296894 70276 297074 70364
rect 297182 70276 297362 70364
rect 297470 70276 297650 70364
rect 297758 70276 297938 70364
rect 298046 70276 298226 70364
rect 298334 70276 298514 70364
rect 310814 70276 310994 70364
rect 311102 70276 311282 70364
rect 311390 70276 311570 70364
rect 311678 70276 311858 70364
rect 311966 70276 312146 70364
rect 312254 70276 312434 70364
rect 312542 70276 312722 70364
rect 312830 70276 313010 70364
rect 325310 70276 325490 70364
rect 325598 70276 325778 70364
rect 325886 70276 326066 70364
rect 326174 70276 326354 70364
rect 326462 70276 326642 70364
rect 326750 70276 326930 70364
rect 327038 70276 327218 70364
rect 327326 70276 327506 70364
rect 339806 70276 339986 70364
rect 340094 70276 340274 70364
rect 340382 70276 340562 70364
rect 340670 70276 340850 70364
rect 340958 70276 341138 70364
rect 341246 70276 341426 70364
rect 341534 70276 341714 70364
rect 341822 70276 342002 70364
rect 354302 70276 354482 70364
rect 354590 70276 354770 70364
rect 354878 70276 355058 70364
rect 355166 70276 355346 70364
rect 355454 70276 355634 70364
rect 355742 70276 355922 70364
rect 356030 70276 356210 70364
rect 356318 70276 356498 70364
rect 368798 70276 368978 70364
rect 369086 70276 369266 70364
rect 369374 70276 369554 70364
rect 369662 70276 369842 70364
rect 369950 70276 370130 70364
rect 370238 70276 370418 70364
rect 370526 70276 370706 70364
rect 370814 70276 370994 70364
rect 383294 70276 383474 70364
rect 383582 70276 383762 70364
rect 383870 70276 384050 70364
rect 384158 70276 384338 70364
rect 384446 70276 384626 70364
rect 384734 70276 384914 70364
rect 385022 70276 385202 70364
rect 385310 70276 385490 70364
rect 397790 70276 397970 70364
rect 398078 70276 398258 70364
rect 398366 70276 398546 70364
rect 398654 70276 398834 70364
rect 398942 70276 399122 70364
rect 399230 70276 399410 70364
rect 399518 70276 399698 70364
rect 399806 70276 399986 70364
rect 412286 70276 412466 70364
rect 412574 70276 412754 70364
rect 412862 70276 413042 70364
rect 413150 70276 413330 70364
rect 413438 70276 413618 70364
rect 413726 70276 413906 70364
rect 414014 70276 414194 70364
rect 414302 70276 414482 70364
rect 426782 70276 426962 70364
rect 427070 70276 427250 70364
rect 427358 70276 427538 70364
rect 427646 70276 427826 70364
rect 427934 70276 428114 70364
rect 428222 70276 428402 70364
rect 428510 70276 428690 70364
rect 428798 70276 428978 70364
rect 441278 70276 441458 70364
rect 441566 70276 441746 70364
rect 441854 70276 442034 70364
rect 442142 70276 442322 70364
rect 442430 70276 442610 70364
rect 442718 70276 442898 70364
rect 443006 70276 443186 70364
rect 443294 70276 443474 70364
rect 455774 70276 455954 70364
rect 456062 70276 456242 70364
rect 456350 70276 456530 70364
rect 456638 70276 456818 70364
rect 456926 70276 457106 70364
rect 457214 70276 457394 70364
rect 457502 70276 457682 70364
rect 457790 70276 457970 70364
rect 180350 70060 180530 70148
rect 180638 70060 180818 70148
rect 180926 70060 181106 70148
rect 181214 70060 181394 70148
rect 181502 70060 181682 70148
rect 181790 70060 181970 70148
rect 182078 70060 182258 70148
rect 182366 70060 182546 70148
rect 194846 70060 195026 70148
rect 195134 70060 195314 70148
rect 195422 70060 195602 70148
rect 195710 70060 195890 70148
rect 195998 70060 196178 70148
rect 196286 70060 196466 70148
rect 196574 70060 196754 70148
rect 196862 70060 197042 70148
rect 209342 70060 209522 70148
rect 209630 70060 209810 70148
rect 209918 70060 210098 70148
rect 210206 70060 210386 70148
rect 210494 70060 210674 70148
rect 210782 70060 210962 70148
rect 211070 70060 211250 70148
rect 211358 70060 211538 70148
rect 223838 70060 224018 70148
rect 224126 70060 224306 70148
rect 224414 70060 224594 70148
rect 224702 70060 224882 70148
rect 224990 70060 225170 70148
rect 225278 70060 225458 70148
rect 225566 70060 225746 70148
rect 225854 70060 226034 70148
rect 238334 70060 238514 70148
rect 238622 70060 238802 70148
rect 238910 70060 239090 70148
rect 239198 70060 239378 70148
rect 239486 70060 239666 70148
rect 239774 70060 239954 70148
rect 240062 70060 240242 70148
rect 240350 70060 240530 70148
rect 252830 70060 253010 70148
rect 253118 70060 253298 70148
rect 253406 70060 253586 70148
rect 253694 70060 253874 70148
rect 253982 70060 254162 70148
rect 254270 70060 254450 70148
rect 254558 70060 254738 70148
rect 254846 70060 255026 70148
rect 267326 70060 267506 70148
rect 267614 70060 267794 70148
rect 267902 70060 268082 70148
rect 268190 70060 268370 70148
rect 268478 70060 268658 70148
rect 268766 70060 268946 70148
rect 269054 70060 269234 70148
rect 269342 70060 269522 70148
rect 281822 70060 282002 70148
rect 282110 70060 282290 70148
rect 282398 70060 282578 70148
rect 282686 70060 282866 70148
rect 282974 70060 283154 70148
rect 283262 70060 283442 70148
rect 283550 70060 283730 70148
rect 283838 70060 284018 70148
rect 296318 70060 296498 70148
rect 296606 70060 296786 70148
rect 296894 70060 297074 70148
rect 297182 70060 297362 70148
rect 297470 70060 297650 70148
rect 297758 70060 297938 70148
rect 298046 70060 298226 70148
rect 298334 70060 298514 70148
rect 310814 70060 310994 70148
rect 311102 70060 311282 70148
rect 311390 70060 311570 70148
rect 311678 70060 311858 70148
rect 311966 70060 312146 70148
rect 312254 70060 312434 70148
rect 312542 70060 312722 70148
rect 312830 70060 313010 70148
rect 325310 70060 325490 70148
rect 325598 70060 325778 70148
rect 325886 70060 326066 70148
rect 326174 70060 326354 70148
rect 326462 70060 326642 70148
rect 326750 70060 326930 70148
rect 327038 70060 327218 70148
rect 327326 70060 327506 70148
rect 339806 70060 339986 70148
rect 340094 70060 340274 70148
rect 340382 70060 340562 70148
rect 340670 70060 340850 70148
rect 340958 70060 341138 70148
rect 341246 70060 341426 70148
rect 341534 70060 341714 70148
rect 341822 70060 342002 70148
rect 354302 70060 354482 70148
rect 354590 70060 354770 70148
rect 354878 70060 355058 70148
rect 355166 70060 355346 70148
rect 355454 70060 355634 70148
rect 355742 70060 355922 70148
rect 356030 70060 356210 70148
rect 356318 70060 356498 70148
rect 368798 70060 368978 70148
rect 369086 70060 369266 70148
rect 369374 70060 369554 70148
rect 369662 70060 369842 70148
rect 369950 70060 370130 70148
rect 370238 70060 370418 70148
rect 370526 70060 370706 70148
rect 370814 70060 370994 70148
rect 383294 70060 383474 70148
rect 383582 70060 383762 70148
rect 383870 70060 384050 70148
rect 384158 70060 384338 70148
rect 384446 70060 384626 70148
rect 384734 70060 384914 70148
rect 385022 70060 385202 70148
rect 385310 70060 385490 70148
rect 397790 70060 397970 70148
rect 398078 70060 398258 70148
rect 398366 70060 398546 70148
rect 398654 70060 398834 70148
rect 398942 70060 399122 70148
rect 399230 70060 399410 70148
rect 399518 70060 399698 70148
rect 399806 70060 399986 70148
rect 412286 70060 412466 70148
rect 412574 70060 412754 70148
rect 412862 70060 413042 70148
rect 413150 70060 413330 70148
rect 413438 70060 413618 70148
rect 413726 70060 413906 70148
rect 414014 70060 414194 70148
rect 414302 70060 414482 70148
rect 426782 70060 426962 70148
rect 427070 70060 427250 70148
rect 427358 70060 427538 70148
rect 427646 70060 427826 70148
rect 427934 70060 428114 70148
rect 428222 70060 428402 70148
rect 428510 70060 428690 70148
rect 428798 70060 428978 70148
rect 441278 70060 441458 70148
rect 441566 70060 441746 70148
rect 441854 70060 442034 70148
rect 442142 70060 442322 70148
rect 442430 70060 442610 70148
rect 442718 70060 442898 70148
rect 443006 70060 443186 70148
rect 443294 70060 443474 70148
rect 455774 70060 455954 70148
rect 456062 70060 456242 70148
rect 456350 70060 456530 70148
rect 456638 70060 456818 70148
rect 456926 70060 457106 70148
rect 457214 70060 457394 70148
rect 457502 70060 457682 70148
rect 457790 70060 457970 70148
rect 180350 55908 180530 55996
rect 180638 55908 180818 55996
rect 180926 55908 181106 55996
rect 181214 55908 181394 55996
rect 181502 55908 181682 55996
rect 181790 55908 181970 55996
rect 182078 55908 182258 55996
rect 182366 55908 182546 55996
rect 194846 55908 195026 55996
rect 195134 55908 195314 55996
rect 195422 55908 195602 55996
rect 195710 55908 195890 55996
rect 195998 55908 196178 55996
rect 196286 55908 196466 55996
rect 196574 55908 196754 55996
rect 196862 55908 197042 55996
rect 209342 55908 209522 55996
rect 209630 55908 209810 55996
rect 209918 55908 210098 55996
rect 210206 55908 210386 55996
rect 210494 55908 210674 55996
rect 210782 55908 210962 55996
rect 211070 55908 211250 55996
rect 211358 55908 211538 55996
rect 223838 55908 224018 55996
rect 224126 55908 224306 55996
rect 224414 55908 224594 55996
rect 224702 55908 224882 55996
rect 224990 55908 225170 55996
rect 225278 55908 225458 55996
rect 225566 55908 225746 55996
rect 225854 55908 226034 55996
rect 238334 55908 238514 55996
rect 238622 55908 238802 55996
rect 238910 55908 239090 55996
rect 239198 55908 239378 55996
rect 239486 55908 239666 55996
rect 239774 55908 239954 55996
rect 240062 55908 240242 55996
rect 240350 55908 240530 55996
rect 252830 55908 253010 55996
rect 253118 55908 253298 55996
rect 253406 55908 253586 55996
rect 253694 55908 253874 55996
rect 253982 55908 254162 55996
rect 254270 55908 254450 55996
rect 254558 55908 254738 55996
rect 254846 55908 255026 55996
rect 267326 55908 267506 55996
rect 267614 55908 267794 55996
rect 267902 55908 268082 55996
rect 268190 55908 268370 55996
rect 268478 55908 268658 55996
rect 268766 55908 268946 55996
rect 269054 55908 269234 55996
rect 269342 55908 269522 55996
rect 281822 55908 282002 55996
rect 282110 55908 282290 55996
rect 282398 55908 282578 55996
rect 282686 55908 282866 55996
rect 282974 55908 283154 55996
rect 283262 55908 283442 55996
rect 283550 55908 283730 55996
rect 283838 55908 284018 55996
rect 296318 55908 296498 55996
rect 296606 55908 296786 55996
rect 296894 55908 297074 55996
rect 297182 55908 297362 55996
rect 297470 55908 297650 55996
rect 297758 55908 297938 55996
rect 298046 55908 298226 55996
rect 298334 55908 298514 55996
rect 310814 55908 310994 55996
rect 311102 55908 311282 55996
rect 311390 55908 311570 55996
rect 311678 55908 311858 55996
rect 311966 55908 312146 55996
rect 312254 55908 312434 55996
rect 312542 55908 312722 55996
rect 312830 55908 313010 55996
rect 325310 55908 325490 55996
rect 325598 55908 325778 55996
rect 325886 55908 326066 55996
rect 326174 55908 326354 55996
rect 326462 55908 326642 55996
rect 326750 55908 326930 55996
rect 327038 55908 327218 55996
rect 327326 55908 327506 55996
rect 339806 55908 339986 55996
rect 340094 55908 340274 55996
rect 340382 55908 340562 55996
rect 340670 55908 340850 55996
rect 340958 55908 341138 55996
rect 341246 55908 341426 55996
rect 341534 55908 341714 55996
rect 341822 55908 342002 55996
rect 354302 55908 354482 55996
rect 354590 55908 354770 55996
rect 354878 55908 355058 55996
rect 355166 55908 355346 55996
rect 355454 55908 355634 55996
rect 355742 55908 355922 55996
rect 356030 55908 356210 55996
rect 356318 55908 356498 55996
rect 368798 55908 368978 55996
rect 369086 55908 369266 55996
rect 369374 55908 369554 55996
rect 369662 55908 369842 55996
rect 369950 55908 370130 55996
rect 370238 55908 370418 55996
rect 370526 55908 370706 55996
rect 370814 55908 370994 55996
rect 383294 55908 383474 55996
rect 383582 55908 383762 55996
rect 383870 55908 384050 55996
rect 384158 55908 384338 55996
rect 384446 55908 384626 55996
rect 384734 55908 384914 55996
rect 385022 55908 385202 55996
rect 385310 55908 385490 55996
rect 397790 55908 397970 55996
rect 398078 55908 398258 55996
rect 398366 55908 398546 55996
rect 398654 55908 398834 55996
rect 398942 55908 399122 55996
rect 399230 55908 399410 55996
rect 399518 55908 399698 55996
rect 399806 55908 399986 55996
rect 412286 55908 412466 55996
rect 412574 55908 412754 55996
rect 412862 55908 413042 55996
rect 413150 55908 413330 55996
rect 413438 55908 413618 55996
rect 413726 55908 413906 55996
rect 414014 55908 414194 55996
rect 414302 55908 414482 55996
rect 426782 55908 426962 55996
rect 427070 55908 427250 55996
rect 427358 55908 427538 55996
rect 427646 55908 427826 55996
rect 427934 55908 428114 55996
rect 428222 55908 428402 55996
rect 428510 55908 428690 55996
rect 428798 55908 428978 55996
rect 441278 55908 441458 55996
rect 441566 55908 441746 55996
rect 441854 55908 442034 55996
rect 442142 55908 442322 55996
rect 442430 55908 442610 55996
rect 442718 55908 442898 55996
rect 443006 55908 443186 55996
rect 443294 55908 443474 55996
rect 455774 55908 455954 55996
rect 456062 55908 456242 55996
rect 456350 55908 456530 55996
rect 456638 55908 456818 55996
rect 456926 55908 457106 55996
rect 457214 55908 457394 55996
rect 457502 55908 457682 55996
rect 457790 55908 457970 55996
rect 180350 55692 180530 55780
rect 180638 55692 180818 55780
rect 180926 55692 181106 55780
rect 181214 55692 181394 55780
rect 181502 55692 181682 55780
rect 181790 55692 181970 55780
rect 182078 55692 182258 55780
rect 182366 55692 182546 55780
rect 194846 55692 195026 55780
rect 195134 55692 195314 55780
rect 195422 55692 195602 55780
rect 195710 55692 195890 55780
rect 195998 55692 196178 55780
rect 196286 55692 196466 55780
rect 196574 55692 196754 55780
rect 196862 55692 197042 55780
rect 209342 55692 209522 55780
rect 209630 55692 209810 55780
rect 209918 55692 210098 55780
rect 210206 55692 210386 55780
rect 210494 55692 210674 55780
rect 210782 55692 210962 55780
rect 211070 55692 211250 55780
rect 211358 55692 211538 55780
rect 223838 55692 224018 55780
rect 224126 55692 224306 55780
rect 224414 55692 224594 55780
rect 224702 55692 224882 55780
rect 224990 55692 225170 55780
rect 225278 55692 225458 55780
rect 225566 55692 225746 55780
rect 225854 55692 226034 55780
rect 238334 55692 238514 55780
rect 238622 55692 238802 55780
rect 238910 55692 239090 55780
rect 239198 55692 239378 55780
rect 239486 55692 239666 55780
rect 239774 55692 239954 55780
rect 240062 55692 240242 55780
rect 240350 55692 240530 55780
rect 252830 55692 253010 55780
rect 253118 55692 253298 55780
rect 253406 55692 253586 55780
rect 253694 55692 253874 55780
rect 253982 55692 254162 55780
rect 254270 55692 254450 55780
rect 254558 55692 254738 55780
rect 254846 55692 255026 55780
rect 267326 55692 267506 55780
rect 267614 55692 267794 55780
rect 267902 55692 268082 55780
rect 268190 55692 268370 55780
rect 268478 55692 268658 55780
rect 268766 55692 268946 55780
rect 269054 55692 269234 55780
rect 269342 55692 269522 55780
rect 281822 55692 282002 55780
rect 282110 55692 282290 55780
rect 282398 55692 282578 55780
rect 282686 55692 282866 55780
rect 282974 55692 283154 55780
rect 283262 55692 283442 55780
rect 283550 55692 283730 55780
rect 283838 55692 284018 55780
rect 296318 55692 296498 55780
rect 296606 55692 296786 55780
rect 296894 55692 297074 55780
rect 297182 55692 297362 55780
rect 297470 55692 297650 55780
rect 297758 55692 297938 55780
rect 298046 55692 298226 55780
rect 298334 55692 298514 55780
rect 310814 55692 310994 55780
rect 311102 55692 311282 55780
rect 311390 55692 311570 55780
rect 311678 55692 311858 55780
rect 311966 55692 312146 55780
rect 312254 55692 312434 55780
rect 312542 55692 312722 55780
rect 312830 55692 313010 55780
rect 325310 55692 325490 55780
rect 325598 55692 325778 55780
rect 325886 55692 326066 55780
rect 326174 55692 326354 55780
rect 326462 55692 326642 55780
rect 326750 55692 326930 55780
rect 327038 55692 327218 55780
rect 327326 55692 327506 55780
rect 339806 55692 339986 55780
rect 340094 55692 340274 55780
rect 340382 55692 340562 55780
rect 340670 55692 340850 55780
rect 340958 55692 341138 55780
rect 341246 55692 341426 55780
rect 341534 55692 341714 55780
rect 341822 55692 342002 55780
rect 354302 55692 354482 55780
rect 354590 55692 354770 55780
rect 354878 55692 355058 55780
rect 355166 55692 355346 55780
rect 355454 55692 355634 55780
rect 355742 55692 355922 55780
rect 356030 55692 356210 55780
rect 356318 55692 356498 55780
rect 368798 55692 368978 55780
rect 369086 55692 369266 55780
rect 369374 55692 369554 55780
rect 369662 55692 369842 55780
rect 369950 55692 370130 55780
rect 370238 55692 370418 55780
rect 370526 55692 370706 55780
rect 370814 55692 370994 55780
rect 383294 55692 383474 55780
rect 383582 55692 383762 55780
rect 383870 55692 384050 55780
rect 384158 55692 384338 55780
rect 384446 55692 384626 55780
rect 384734 55692 384914 55780
rect 385022 55692 385202 55780
rect 385310 55692 385490 55780
rect 397790 55692 397970 55780
rect 398078 55692 398258 55780
rect 398366 55692 398546 55780
rect 398654 55692 398834 55780
rect 398942 55692 399122 55780
rect 399230 55692 399410 55780
rect 399518 55692 399698 55780
rect 399806 55692 399986 55780
rect 412286 55692 412466 55780
rect 412574 55692 412754 55780
rect 412862 55692 413042 55780
rect 413150 55692 413330 55780
rect 413438 55692 413618 55780
rect 413726 55692 413906 55780
rect 414014 55692 414194 55780
rect 414302 55692 414482 55780
rect 426782 55692 426962 55780
rect 427070 55692 427250 55780
rect 427358 55692 427538 55780
rect 427646 55692 427826 55780
rect 427934 55692 428114 55780
rect 428222 55692 428402 55780
rect 428510 55692 428690 55780
rect 428798 55692 428978 55780
rect 441278 55692 441458 55780
rect 441566 55692 441746 55780
rect 441854 55692 442034 55780
rect 442142 55692 442322 55780
rect 442430 55692 442610 55780
rect 442718 55692 442898 55780
rect 443006 55692 443186 55780
rect 443294 55692 443474 55780
rect 455774 55692 455954 55780
rect 456062 55692 456242 55780
rect 456350 55692 456530 55780
rect 456638 55692 456818 55780
rect 456926 55692 457106 55780
rect 457214 55692 457394 55780
rect 457502 55692 457682 55780
rect 457790 55692 457970 55780
rect 180350 55216 180530 55304
rect 180638 55216 180818 55304
rect 180926 55216 181106 55304
rect 181214 55216 181394 55304
rect 181502 55216 181682 55304
rect 181790 55216 181970 55304
rect 182078 55216 182258 55304
rect 182366 55216 182546 55304
rect 194846 55216 195026 55304
rect 195134 55216 195314 55304
rect 195422 55216 195602 55304
rect 195710 55216 195890 55304
rect 195998 55216 196178 55304
rect 196286 55216 196466 55304
rect 196574 55216 196754 55304
rect 196862 55216 197042 55304
rect 209342 55216 209522 55304
rect 209630 55216 209810 55304
rect 209918 55216 210098 55304
rect 210206 55216 210386 55304
rect 210494 55216 210674 55304
rect 210782 55216 210962 55304
rect 211070 55216 211250 55304
rect 211358 55216 211538 55304
rect 223838 55216 224018 55304
rect 224126 55216 224306 55304
rect 224414 55216 224594 55304
rect 224702 55216 224882 55304
rect 224990 55216 225170 55304
rect 225278 55216 225458 55304
rect 225566 55216 225746 55304
rect 225854 55216 226034 55304
rect 238334 55216 238514 55304
rect 238622 55216 238802 55304
rect 238910 55216 239090 55304
rect 239198 55216 239378 55304
rect 239486 55216 239666 55304
rect 239774 55216 239954 55304
rect 240062 55216 240242 55304
rect 240350 55216 240530 55304
rect 252830 55216 253010 55304
rect 253118 55216 253298 55304
rect 253406 55216 253586 55304
rect 253694 55216 253874 55304
rect 253982 55216 254162 55304
rect 254270 55216 254450 55304
rect 254558 55216 254738 55304
rect 254846 55216 255026 55304
rect 267326 55216 267506 55304
rect 267614 55216 267794 55304
rect 267902 55216 268082 55304
rect 268190 55216 268370 55304
rect 268478 55216 268658 55304
rect 268766 55216 268946 55304
rect 269054 55216 269234 55304
rect 269342 55216 269522 55304
rect 281822 55216 282002 55304
rect 282110 55216 282290 55304
rect 282398 55216 282578 55304
rect 282686 55216 282866 55304
rect 282974 55216 283154 55304
rect 283262 55216 283442 55304
rect 283550 55216 283730 55304
rect 283838 55216 284018 55304
rect 296318 55216 296498 55304
rect 296606 55216 296786 55304
rect 296894 55216 297074 55304
rect 297182 55216 297362 55304
rect 297470 55216 297650 55304
rect 297758 55216 297938 55304
rect 298046 55216 298226 55304
rect 298334 55216 298514 55304
rect 310814 55216 310994 55304
rect 311102 55216 311282 55304
rect 311390 55216 311570 55304
rect 311678 55216 311858 55304
rect 311966 55216 312146 55304
rect 312254 55216 312434 55304
rect 312542 55216 312722 55304
rect 312830 55216 313010 55304
rect 325310 55216 325490 55304
rect 325598 55216 325778 55304
rect 325886 55216 326066 55304
rect 326174 55216 326354 55304
rect 326462 55216 326642 55304
rect 326750 55216 326930 55304
rect 327038 55216 327218 55304
rect 327326 55216 327506 55304
rect 339806 55216 339986 55304
rect 340094 55216 340274 55304
rect 340382 55216 340562 55304
rect 340670 55216 340850 55304
rect 340958 55216 341138 55304
rect 341246 55216 341426 55304
rect 341534 55216 341714 55304
rect 341822 55216 342002 55304
rect 354302 55216 354482 55304
rect 354590 55216 354770 55304
rect 354878 55216 355058 55304
rect 355166 55216 355346 55304
rect 355454 55216 355634 55304
rect 355742 55216 355922 55304
rect 356030 55216 356210 55304
rect 356318 55216 356498 55304
rect 368798 55216 368978 55304
rect 369086 55216 369266 55304
rect 369374 55216 369554 55304
rect 369662 55216 369842 55304
rect 369950 55216 370130 55304
rect 370238 55216 370418 55304
rect 370526 55216 370706 55304
rect 370814 55216 370994 55304
rect 383294 55216 383474 55304
rect 383582 55216 383762 55304
rect 383870 55216 384050 55304
rect 384158 55216 384338 55304
rect 384446 55216 384626 55304
rect 384734 55216 384914 55304
rect 385022 55216 385202 55304
rect 385310 55216 385490 55304
rect 397790 55216 397970 55304
rect 398078 55216 398258 55304
rect 398366 55216 398546 55304
rect 398654 55216 398834 55304
rect 398942 55216 399122 55304
rect 399230 55216 399410 55304
rect 399518 55216 399698 55304
rect 399806 55216 399986 55304
rect 412286 55216 412466 55304
rect 412574 55216 412754 55304
rect 412862 55216 413042 55304
rect 413150 55216 413330 55304
rect 413438 55216 413618 55304
rect 413726 55216 413906 55304
rect 414014 55216 414194 55304
rect 414302 55216 414482 55304
rect 426782 55216 426962 55304
rect 427070 55216 427250 55304
rect 427358 55216 427538 55304
rect 427646 55216 427826 55304
rect 427934 55216 428114 55304
rect 428222 55216 428402 55304
rect 428510 55216 428690 55304
rect 428798 55216 428978 55304
rect 441278 55216 441458 55304
rect 441566 55216 441746 55304
rect 441854 55216 442034 55304
rect 442142 55216 442322 55304
rect 442430 55216 442610 55304
rect 442718 55216 442898 55304
rect 443006 55216 443186 55304
rect 443294 55216 443474 55304
rect 455774 55216 455954 55304
rect 456062 55216 456242 55304
rect 456350 55216 456530 55304
rect 456638 55216 456818 55304
rect 456926 55216 457106 55304
rect 457214 55216 457394 55304
rect 457502 55216 457682 55304
rect 457790 55216 457970 55304
rect 180350 55000 180530 55088
rect 180638 55000 180818 55088
rect 180926 55000 181106 55088
rect 181214 55000 181394 55088
rect 181502 55000 181682 55088
rect 181790 55000 181970 55088
rect 182078 55000 182258 55088
rect 182366 55000 182546 55088
rect 194846 55000 195026 55088
rect 195134 55000 195314 55088
rect 195422 55000 195602 55088
rect 195710 55000 195890 55088
rect 195998 55000 196178 55088
rect 196286 55000 196466 55088
rect 196574 55000 196754 55088
rect 196862 55000 197042 55088
rect 209342 55000 209522 55088
rect 209630 55000 209810 55088
rect 209918 55000 210098 55088
rect 210206 55000 210386 55088
rect 210494 55000 210674 55088
rect 210782 55000 210962 55088
rect 211070 55000 211250 55088
rect 211358 55000 211538 55088
rect 223838 55000 224018 55088
rect 224126 55000 224306 55088
rect 224414 55000 224594 55088
rect 224702 55000 224882 55088
rect 224990 55000 225170 55088
rect 225278 55000 225458 55088
rect 225566 55000 225746 55088
rect 225854 55000 226034 55088
rect 238334 55000 238514 55088
rect 238622 55000 238802 55088
rect 238910 55000 239090 55088
rect 239198 55000 239378 55088
rect 239486 55000 239666 55088
rect 239774 55000 239954 55088
rect 240062 55000 240242 55088
rect 240350 55000 240530 55088
rect 252830 55000 253010 55088
rect 253118 55000 253298 55088
rect 253406 55000 253586 55088
rect 253694 55000 253874 55088
rect 253982 55000 254162 55088
rect 254270 55000 254450 55088
rect 254558 55000 254738 55088
rect 254846 55000 255026 55088
rect 267326 55000 267506 55088
rect 267614 55000 267794 55088
rect 267902 55000 268082 55088
rect 268190 55000 268370 55088
rect 268478 55000 268658 55088
rect 268766 55000 268946 55088
rect 269054 55000 269234 55088
rect 269342 55000 269522 55088
rect 281822 55000 282002 55088
rect 282110 55000 282290 55088
rect 282398 55000 282578 55088
rect 282686 55000 282866 55088
rect 282974 55000 283154 55088
rect 283262 55000 283442 55088
rect 283550 55000 283730 55088
rect 283838 55000 284018 55088
rect 296318 55000 296498 55088
rect 296606 55000 296786 55088
rect 296894 55000 297074 55088
rect 297182 55000 297362 55088
rect 297470 55000 297650 55088
rect 297758 55000 297938 55088
rect 298046 55000 298226 55088
rect 298334 55000 298514 55088
rect 310814 55000 310994 55088
rect 311102 55000 311282 55088
rect 311390 55000 311570 55088
rect 311678 55000 311858 55088
rect 311966 55000 312146 55088
rect 312254 55000 312434 55088
rect 312542 55000 312722 55088
rect 312830 55000 313010 55088
rect 325310 55000 325490 55088
rect 325598 55000 325778 55088
rect 325886 55000 326066 55088
rect 326174 55000 326354 55088
rect 326462 55000 326642 55088
rect 326750 55000 326930 55088
rect 327038 55000 327218 55088
rect 327326 55000 327506 55088
rect 339806 55000 339986 55088
rect 340094 55000 340274 55088
rect 340382 55000 340562 55088
rect 340670 55000 340850 55088
rect 340958 55000 341138 55088
rect 341246 55000 341426 55088
rect 341534 55000 341714 55088
rect 341822 55000 342002 55088
rect 354302 55000 354482 55088
rect 354590 55000 354770 55088
rect 354878 55000 355058 55088
rect 355166 55000 355346 55088
rect 355454 55000 355634 55088
rect 355742 55000 355922 55088
rect 356030 55000 356210 55088
rect 356318 55000 356498 55088
rect 368798 55000 368978 55088
rect 369086 55000 369266 55088
rect 369374 55000 369554 55088
rect 369662 55000 369842 55088
rect 369950 55000 370130 55088
rect 370238 55000 370418 55088
rect 370526 55000 370706 55088
rect 370814 55000 370994 55088
rect 383294 55000 383474 55088
rect 383582 55000 383762 55088
rect 383870 55000 384050 55088
rect 384158 55000 384338 55088
rect 384446 55000 384626 55088
rect 384734 55000 384914 55088
rect 385022 55000 385202 55088
rect 385310 55000 385490 55088
rect 397790 55000 397970 55088
rect 398078 55000 398258 55088
rect 398366 55000 398546 55088
rect 398654 55000 398834 55088
rect 398942 55000 399122 55088
rect 399230 55000 399410 55088
rect 399518 55000 399698 55088
rect 399806 55000 399986 55088
rect 412286 55000 412466 55088
rect 412574 55000 412754 55088
rect 412862 55000 413042 55088
rect 413150 55000 413330 55088
rect 413438 55000 413618 55088
rect 413726 55000 413906 55088
rect 414014 55000 414194 55088
rect 414302 55000 414482 55088
rect 426782 55000 426962 55088
rect 427070 55000 427250 55088
rect 427358 55000 427538 55088
rect 427646 55000 427826 55088
rect 427934 55000 428114 55088
rect 428222 55000 428402 55088
rect 428510 55000 428690 55088
rect 428798 55000 428978 55088
rect 441278 55000 441458 55088
rect 441566 55000 441746 55088
rect 441854 55000 442034 55088
rect 442142 55000 442322 55088
rect 442430 55000 442610 55088
rect 442718 55000 442898 55088
rect 443006 55000 443186 55088
rect 443294 55000 443474 55088
rect 455774 55000 455954 55088
rect 456062 55000 456242 55088
rect 456350 55000 456530 55088
rect 456638 55000 456818 55088
rect 456926 55000 457106 55088
rect 457214 55000 457394 55088
rect 457502 55000 457682 55088
rect 457790 55000 457970 55088
rect 180350 40848 180530 40936
rect 180638 40848 180818 40936
rect 180926 40848 181106 40936
rect 181214 40848 181394 40936
rect 181502 40848 181682 40936
rect 181790 40848 181970 40936
rect 182078 40848 182258 40936
rect 182366 40848 182546 40936
rect 194846 40848 195026 40936
rect 195134 40848 195314 40936
rect 195422 40848 195602 40936
rect 195710 40848 195890 40936
rect 195998 40848 196178 40936
rect 196286 40848 196466 40936
rect 196574 40848 196754 40936
rect 196862 40848 197042 40936
rect 209342 40848 209522 40936
rect 209630 40848 209810 40936
rect 209918 40848 210098 40936
rect 210206 40848 210386 40936
rect 210494 40848 210674 40936
rect 210782 40848 210962 40936
rect 211070 40848 211250 40936
rect 211358 40848 211538 40936
rect 223838 40848 224018 40936
rect 224126 40848 224306 40936
rect 224414 40848 224594 40936
rect 224702 40848 224882 40936
rect 224990 40848 225170 40936
rect 225278 40848 225458 40936
rect 225566 40848 225746 40936
rect 225854 40848 226034 40936
rect 238334 40848 238514 40936
rect 238622 40848 238802 40936
rect 238910 40848 239090 40936
rect 239198 40848 239378 40936
rect 239486 40848 239666 40936
rect 239774 40848 239954 40936
rect 240062 40848 240242 40936
rect 240350 40848 240530 40936
rect 252830 40848 253010 40936
rect 253118 40848 253298 40936
rect 253406 40848 253586 40936
rect 253694 40848 253874 40936
rect 253982 40848 254162 40936
rect 254270 40848 254450 40936
rect 254558 40848 254738 40936
rect 254846 40848 255026 40936
rect 267326 40848 267506 40936
rect 267614 40848 267794 40936
rect 267902 40848 268082 40936
rect 268190 40848 268370 40936
rect 268478 40848 268658 40936
rect 268766 40848 268946 40936
rect 269054 40848 269234 40936
rect 269342 40848 269522 40936
rect 281822 40848 282002 40936
rect 282110 40848 282290 40936
rect 282398 40848 282578 40936
rect 282686 40848 282866 40936
rect 282974 40848 283154 40936
rect 283262 40848 283442 40936
rect 283550 40848 283730 40936
rect 283838 40848 284018 40936
rect 296318 40848 296498 40936
rect 296606 40848 296786 40936
rect 296894 40848 297074 40936
rect 297182 40848 297362 40936
rect 297470 40848 297650 40936
rect 297758 40848 297938 40936
rect 298046 40848 298226 40936
rect 298334 40848 298514 40936
rect 310814 40848 310994 40936
rect 311102 40848 311282 40936
rect 311390 40848 311570 40936
rect 311678 40848 311858 40936
rect 311966 40848 312146 40936
rect 312254 40848 312434 40936
rect 312542 40848 312722 40936
rect 312830 40848 313010 40936
rect 325310 40848 325490 40936
rect 325598 40848 325778 40936
rect 325886 40848 326066 40936
rect 326174 40848 326354 40936
rect 326462 40848 326642 40936
rect 326750 40848 326930 40936
rect 327038 40848 327218 40936
rect 327326 40848 327506 40936
rect 339806 40848 339986 40936
rect 340094 40848 340274 40936
rect 340382 40848 340562 40936
rect 340670 40848 340850 40936
rect 340958 40848 341138 40936
rect 341246 40848 341426 40936
rect 341534 40848 341714 40936
rect 341822 40848 342002 40936
rect 354302 40848 354482 40936
rect 354590 40848 354770 40936
rect 354878 40848 355058 40936
rect 355166 40848 355346 40936
rect 355454 40848 355634 40936
rect 355742 40848 355922 40936
rect 356030 40848 356210 40936
rect 356318 40848 356498 40936
rect 368798 40848 368978 40936
rect 369086 40848 369266 40936
rect 369374 40848 369554 40936
rect 369662 40848 369842 40936
rect 369950 40848 370130 40936
rect 370238 40848 370418 40936
rect 370526 40848 370706 40936
rect 370814 40848 370994 40936
rect 383294 40848 383474 40936
rect 383582 40848 383762 40936
rect 383870 40848 384050 40936
rect 384158 40848 384338 40936
rect 384446 40848 384626 40936
rect 384734 40848 384914 40936
rect 385022 40848 385202 40936
rect 385310 40848 385490 40936
rect 397790 40848 397970 40936
rect 398078 40848 398258 40936
rect 398366 40848 398546 40936
rect 398654 40848 398834 40936
rect 398942 40848 399122 40936
rect 399230 40848 399410 40936
rect 399518 40848 399698 40936
rect 399806 40848 399986 40936
rect 412286 40848 412466 40936
rect 412574 40848 412754 40936
rect 412862 40848 413042 40936
rect 413150 40848 413330 40936
rect 413438 40848 413618 40936
rect 413726 40848 413906 40936
rect 414014 40848 414194 40936
rect 414302 40848 414482 40936
rect 426782 40848 426962 40936
rect 427070 40848 427250 40936
rect 427358 40848 427538 40936
rect 427646 40848 427826 40936
rect 427934 40848 428114 40936
rect 428222 40848 428402 40936
rect 428510 40848 428690 40936
rect 428798 40848 428978 40936
rect 441278 40848 441458 40936
rect 441566 40848 441746 40936
rect 441854 40848 442034 40936
rect 442142 40848 442322 40936
rect 442430 40848 442610 40936
rect 442718 40848 442898 40936
rect 443006 40848 443186 40936
rect 443294 40848 443474 40936
rect 455774 40848 455954 40936
rect 456062 40848 456242 40936
rect 456350 40848 456530 40936
rect 456638 40848 456818 40936
rect 456926 40848 457106 40936
rect 457214 40848 457394 40936
rect 457502 40848 457682 40936
rect 457790 40848 457970 40936
rect 180350 40632 180530 40720
rect 180638 40632 180818 40720
rect 180926 40632 181106 40720
rect 181214 40632 181394 40720
rect 181502 40632 181682 40720
rect 181790 40632 181970 40720
rect 182078 40632 182258 40720
rect 182366 40632 182546 40720
rect 194846 40632 195026 40720
rect 195134 40632 195314 40720
rect 195422 40632 195602 40720
rect 195710 40632 195890 40720
rect 195998 40632 196178 40720
rect 196286 40632 196466 40720
rect 196574 40632 196754 40720
rect 196862 40632 197042 40720
rect 209342 40632 209522 40720
rect 209630 40632 209810 40720
rect 209918 40632 210098 40720
rect 210206 40632 210386 40720
rect 210494 40632 210674 40720
rect 210782 40632 210962 40720
rect 211070 40632 211250 40720
rect 211358 40632 211538 40720
rect 223838 40632 224018 40720
rect 224126 40632 224306 40720
rect 224414 40632 224594 40720
rect 224702 40632 224882 40720
rect 224990 40632 225170 40720
rect 225278 40632 225458 40720
rect 225566 40632 225746 40720
rect 225854 40632 226034 40720
rect 238334 40632 238514 40720
rect 238622 40632 238802 40720
rect 238910 40632 239090 40720
rect 239198 40632 239378 40720
rect 239486 40632 239666 40720
rect 239774 40632 239954 40720
rect 240062 40632 240242 40720
rect 240350 40632 240530 40720
rect 252830 40632 253010 40720
rect 253118 40632 253298 40720
rect 253406 40632 253586 40720
rect 253694 40632 253874 40720
rect 253982 40632 254162 40720
rect 254270 40632 254450 40720
rect 254558 40632 254738 40720
rect 254846 40632 255026 40720
rect 267326 40632 267506 40720
rect 267614 40632 267794 40720
rect 267902 40632 268082 40720
rect 268190 40632 268370 40720
rect 268478 40632 268658 40720
rect 268766 40632 268946 40720
rect 269054 40632 269234 40720
rect 269342 40632 269522 40720
rect 281822 40632 282002 40720
rect 282110 40632 282290 40720
rect 282398 40632 282578 40720
rect 282686 40632 282866 40720
rect 282974 40632 283154 40720
rect 283262 40632 283442 40720
rect 283550 40632 283730 40720
rect 283838 40632 284018 40720
rect 296318 40632 296498 40720
rect 296606 40632 296786 40720
rect 296894 40632 297074 40720
rect 297182 40632 297362 40720
rect 297470 40632 297650 40720
rect 297758 40632 297938 40720
rect 298046 40632 298226 40720
rect 298334 40632 298514 40720
rect 310814 40632 310994 40720
rect 311102 40632 311282 40720
rect 311390 40632 311570 40720
rect 311678 40632 311858 40720
rect 311966 40632 312146 40720
rect 312254 40632 312434 40720
rect 312542 40632 312722 40720
rect 312830 40632 313010 40720
rect 325310 40632 325490 40720
rect 325598 40632 325778 40720
rect 325886 40632 326066 40720
rect 326174 40632 326354 40720
rect 326462 40632 326642 40720
rect 326750 40632 326930 40720
rect 327038 40632 327218 40720
rect 327326 40632 327506 40720
rect 339806 40632 339986 40720
rect 340094 40632 340274 40720
rect 340382 40632 340562 40720
rect 340670 40632 340850 40720
rect 340958 40632 341138 40720
rect 341246 40632 341426 40720
rect 341534 40632 341714 40720
rect 341822 40632 342002 40720
rect 354302 40632 354482 40720
rect 354590 40632 354770 40720
rect 354878 40632 355058 40720
rect 355166 40632 355346 40720
rect 355454 40632 355634 40720
rect 355742 40632 355922 40720
rect 356030 40632 356210 40720
rect 356318 40632 356498 40720
rect 368798 40632 368978 40720
rect 369086 40632 369266 40720
rect 369374 40632 369554 40720
rect 369662 40632 369842 40720
rect 369950 40632 370130 40720
rect 370238 40632 370418 40720
rect 370526 40632 370706 40720
rect 370814 40632 370994 40720
rect 383294 40632 383474 40720
rect 383582 40632 383762 40720
rect 383870 40632 384050 40720
rect 384158 40632 384338 40720
rect 384446 40632 384626 40720
rect 384734 40632 384914 40720
rect 385022 40632 385202 40720
rect 385310 40632 385490 40720
rect 397790 40632 397970 40720
rect 398078 40632 398258 40720
rect 398366 40632 398546 40720
rect 398654 40632 398834 40720
rect 398942 40632 399122 40720
rect 399230 40632 399410 40720
rect 399518 40632 399698 40720
rect 399806 40632 399986 40720
rect 412286 40632 412466 40720
rect 412574 40632 412754 40720
rect 412862 40632 413042 40720
rect 413150 40632 413330 40720
rect 413438 40632 413618 40720
rect 413726 40632 413906 40720
rect 414014 40632 414194 40720
rect 414302 40632 414482 40720
rect 426782 40632 426962 40720
rect 427070 40632 427250 40720
rect 427358 40632 427538 40720
rect 427646 40632 427826 40720
rect 427934 40632 428114 40720
rect 428222 40632 428402 40720
rect 428510 40632 428690 40720
rect 428798 40632 428978 40720
rect 441278 40632 441458 40720
rect 441566 40632 441746 40720
rect 441854 40632 442034 40720
rect 442142 40632 442322 40720
rect 442430 40632 442610 40720
rect 442718 40632 442898 40720
rect 443006 40632 443186 40720
rect 443294 40632 443474 40720
rect 455774 40632 455954 40720
rect 456062 40632 456242 40720
rect 456350 40632 456530 40720
rect 456638 40632 456818 40720
rect 456926 40632 457106 40720
rect 457214 40632 457394 40720
rect 457502 40632 457682 40720
rect 457790 40632 457970 40720
rect 180350 40156 180530 40244
rect 180638 40156 180818 40244
rect 180926 40156 181106 40244
rect 181214 40156 181394 40244
rect 181502 40156 181682 40244
rect 181790 40156 181970 40244
rect 182078 40156 182258 40244
rect 182366 40156 182546 40244
rect 194846 40156 195026 40244
rect 195134 40156 195314 40244
rect 195422 40156 195602 40244
rect 195710 40156 195890 40244
rect 195998 40156 196178 40244
rect 196286 40156 196466 40244
rect 196574 40156 196754 40244
rect 196862 40156 197042 40244
rect 209342 40156 209522 40244
rect 209630 40156 209810 40244
rect 209918 40156 210098 40244
rect 210206 40156 210386 40244
rect 210494 40156 210674 40244
rect 210782 40156 210962 40244
rect 211070 40156 211250 40244
rect 211358 40156 211538 40244
rect 223838 40156 224018 40244
rect 224126 40156 224306 40244
rect 224414 40156 224594 40244
rect 224702 40156 224882 40244
rect 224990 40156 225170 40244
rect 225278 40156 225458 40244
rect 225566 40156 225746 40244
rect 225854 40156 226034 40244
rect 238334 40156 238514 40244
rect 238622 40156 238802 40244
rect 238910 40156 239090 40244
rect 239198 40156 239378 40244
rect 239486 40156 239666 40244
rect 239774 40156 239954 40244
rect 240062 40156 240242 40244
rect 240350 40156 240530 40244
rect 252830 40156 253010 40244
rect 253118 40156 253298 40244
rect 253406 40156 253586 40244
rect 253694 40156 253874 40244
rect 253982 40156 254162 40244
rect 254270 40156 254450 40244
rect 254558 40156 254738 40244
rect 254846 40156 255026 40244
rect 267326 40156 267506 40244
rect 267614 40156 267794 40244
rect 267902 40156 268082 40244
rect 268190 40156 268370 40244
rect 268478 40156 268658 40244
rect 268766 40156 268946 40244
rect 269054 40156 269234 40244
rect 269342 40156 269522 40244
rect 281822 40156 282002 40244
rect 282110 40156 282290 40244
rect 282398 40156 282578 40244
rect 282686 40156 282866 40244
rect 282974 40156 283154 40244
rect 283262 40156 283442 40244
rect 283550 40156 283730 40244
rect 283838 40156 284018 40244
rect 296318 40156 296498 40244
rect 296606 40156 296786 40244
rect 296894 40156 297074 40244
rect 297182 40156 297362 40244
rect 297470 40156 297650 40244
rect 297758 40156 297938 40244
rect 298046 40156 298226 40244
rect 298334 40156 298514 40244
rect 310814 40156 310994 40244
rect 311102 40156 311282 40244
rect 311390 40156 311570 40244
rect 311678 40156 311858 40244
rect 311966 40156 312146 40244
rect 312254 40156 312434 40244
rect 312542 40156 312722 40244
rect 312830 40156 313010 40244
rect 325310 40156 325490 40244
rect 325598 40156 325778 40244
rect 325886 40156 326066 40244
rect 326174 40156 326354 40244
rect 326462 40156 326642 40244
rect 326750 40156 326930 40244
rect 327038 40156 327218 40244
rect 327326 40156 327506 40244
rect 339806 40156 339986 40244
rect 340094 40156 340274 40244
rect 340382 40156 340562 40244
rect 340670 40156 340850 40244
rect 340958 40156 341138 40244
rect 341246 40156 341426 40244
rect 341534 40156 341714 40244
rect 341822 40156 342002 40244
rect 354302 40156 354482 40244
rect 354590 40156 354770 40244
rect 354878 40156 355058 40244
rect 355166 40156 355346 40244
rect 355454 40156 355634 40244
rect 355742 40156 355922 40244
rect 356030 40156 356210 40244
rect 356318 40156 356498 40244
rect 368798 40156 368978 40244
rect 369086 40156 369266 40244
rect 369374 40156 369554 40244
rect 369662 40156 369842 40244
rect 369950 40156 370130 40244
rect 370238 40156 370418 40244
rect 370526 40156 370706 40244
rect 370814 40156 370994 40244
rect 383294 40156 383474 40244
rect 383582 40156 383762 40244
rect 383870 40156 384050 40244
rect 384158 40156 384338 40244
rect 384446 40156 384626 40244
rect 384734 40156 384914 40244
rect 385022 40156 385202 40244
rect 385310 40156 385490 40244
rect 397790 40156 397970 40244
rect 398078 40156 398258 40244
rect 398366 40156 398546 40244
rect 398654 40156 398834 40244
rect 398942 40156 399122 40244
rect 399230 40156 399410 40244
rect 399518 40156 399698 40244
rect 399806 40156 399986 40244
rect 412286 40156 412466 40244
rect 412574 40156 412754 40244
rect 412862 40156 413042 40244
rect 413150 40156 413330 40244
rect 413438 40156 413618 40244
rect 413726 40156 413906 40244
rect 414014 40156 414194 40244
rect 414302 40156 414482 40244
rect 426782 40156 426962 40244
rect 427070 40156 427250 40244
rect 427358 40156 427538 40244
rect 427646 40156 427826 40244
rect 427934 40156 428114 40244
rect 428222 40156 428402 40244
rect 428510 40156 428690 40244
rect 428798 40156 428978 40244
rect 441278 40156 441458 40244
rect 441566 40156 441746 40244
rect 441854 40156 442034 40244
rect 442142 40156 442322 40244
rect 442430 40156 442610 40244
rect 442718 40156 442898 40244
rect 443006 40156 443186 40244
rect 443294 40156 443474 40244
rect 455774 40156 455954 40244
rect 456062 40156 456242 40244
rect 456350 40156 456530 40244
rect 456638 40156 456818 40244
rect 456926 40156 457106 40244
rect 457214 40156 457394 40244
rect 457502 40156 457682 40244
rect 457790 40156 457970 40244
rect 180350 39940 180530 40028
rect 180638 39940 180818 40028
rect 180926 39940 181106 40028
rect 181214 39940 181394 40028
rect 181502 39940 181682 40028
rect 181790 39940 181970 40028
rect 182078 39940 182258 40028
rect 182366 39940 182546 40028
rect 194846 39940 195026 40028
rect 195134 39940 195314 40028
rect 195422 39940 195602 40028
rect 195710 39940 195890 40028
rect 195998 39940 196178 40028
rect 196286 39940 196466 40028
rect 196574 39940 196754 40028
rect 196862 39940 197042 40028
rect 209342 39940 209522 40028
rect 209630 39940 209810 40028
rect 209918 39940 210098 40028
rect 210206 39940 210386 40028
rect 210494 39940 210674 40028
rect 210782 39940 210962 40028
rect 211070 39940 211250 40028
rect 211358 39940 211538 40028
rect 223838 39940 224018 40028
rect 224126 39940 224306 40028
rect 224414 39940 224594 40028
rect 224702 39940 224882 40028
rect 224990 39940 225170 40028
rect 225278 39940 225458 40028
rect 225566 39940 225746 40028
rect 225854 39940 226034 40028
rect 238334 39940 238514 40028
rect 238622 39940 238802 40028
rect 238910 39940 239090 40028
rect 239198 39940 239378 40028
rect 239486 39940 239666 40028
rect 239774 39940 239954 40028
rect 240062 39940 240242 40028
rect 240350 39940 240530 40028
rect 252830 39940 253010 40028
rect 253118 39940 253298 40028
rect 253406 39940 253586 40028
rect 253694 39940 253874 40028
rect 253982 39940 254162 40028
rect 254270 39940 254450 40028
rect 254558 39940 254738 40028
rect 254846 39940 255026 40028
rect 267326 39940 267506 40028
rect 267614 39940 267794 40028
rect 267902 39940 268082 40028
rect 268190 39940 268370 40028
rect 268478 39940 268658 40028
rect 268766 39940 268946 40028
rect 269054 39940 269234 40028
rect 269342 39940 269522 40028
rect 281822 39940 282002 40028
rect 282110 39940 282290 40028
rect 282398 39940 282578 40028
rect 282686 39940 282866 40028
rect 282974 39940 283154 40028
rect 283262 39940 283442 40028
rect 283550 39940 283730 40028
rect 283838 39940 284018 40028
rect 296318 39940 296498 40028
rect 296606 39940 296786 40028
rect 296894 39940 297074 40028
rect 297182 39940 297362 40028
rect 297470 39940 297650 40028
rect 297758 39940 297938 40028
rect 298046 39940 298226 40028
rect 298334 39940 298514 40028
rect 310814 39940 310994 40028
rect 311102 39940 311282 40028
rect 311390 39940 311570 40028
rect 311678 39940 311858 40028
rect 311966 39940 312146 40028
rect 312254 39940 312434 40028
rect 312542 39940 312722 40028
rect 312830 39940 313010 40028
rect 325310 39940 325490 40028
rect 325598 39940 325778 40028
rect 325886 39940 326066 40028
rect 326174 39940 326354 40028
rect 326462 39940 326642 40028
rect 326750 39940 326930 40028
rect 327038 39940 327218 40028
rect 327326 39940 327506 40028
rect 339806 39940 339986 40028
rect 340094 39940 340274 40028
rect 340382 39940 340562 40028
rect 340670 39940 340850 40028
rect 340958 39940 341138 40028
rect 341246 39940 341426 40028
rect 341534 39940 341714 40028
rect 341822 39940 342002 40028
rect 354302 39940 354482 40028
rect 354590 39940 354770 40028
rect 354878 39940 355058 40028
rect 355166 39940 355346 40028
rect 355454 39940 355634 40028
rect 355742 39940 355922 40028
rect 356030 39940 356210 40028
rect 356318 39940 356498 40028
rect 368798 39940 368978 40028
rect 369086 39940 369266 40028
rect 369374 39940 369554 40028
rect 369662 39940 369842 40028
rect 369950 39940 370130 40028
rect 370238 39940 370418 40028
rect 370526 39940 370706 40028
rect 370814 39940 370994 40028
rect 383294 39940 383474 40028
rect 383582 39940 383762 40028
rect 383870 39940 384050 40028
rect 384158 39940 384338 40028
rect 384446 39940 384626 40028
rect 384734 39940 384914 40028
rect 385022 39940 385202 40028
rect 385310 39940 385490 40028
rect 397790 39940 397970 40028
rect 398078 39940 398258 40028
rect 398366 39940 398546 40028
rect 398654 39940 398834 40028
rect 398942 39940 399122 40028
rect 399230 39940 399410 40028
rect 399518 39940 399698 40028
rect 399806 39940 399986 40028
rect 412286 39940 412466 40028
rect 412574 39940 412754 40028
rect 412862 39940 413042 40028
rect 413150 39940 413330 40028
rect 413438 39940 413618 40028
rect 413726 39940 413906 40028
rect 414014 39940 414194 40028
rect 414302 39940 414482 40028
rect 426782 39940 426962 40028
rect 427070 39940 427250 40028
rect 427358 39940 427538 40028
rect 427646 39940 427826 40028
rect 427934 39940 428114 40028
rect 428222 39940 428402 40028
rect 428510 39940 428690 40028
rect 428798 39940 428978 40028
rect 441278 39940 441458 40028
rect 441566 39940 441746 40028
rect 441854 39940 442034 40028
rect 442142 39940 442322 40028
rect 442430 39940 442610 40028
rect 442718 39940 442898 40028
rect 443006 39940 443186 40028
rect 443294 39940 443474 40028
rect 455774 39940 455954 40028
rect 456062 39940 456242 40028
rect 456350 39940 456530 40028
rect 456638 39940 456818 40028
rect 456926 39940 457106 40028
rect 457214 39940 457394 40028
rect 457502 39940 457682 40028
rect 457790 39940 457970 40028
<< dnwell >>
rect 21184 30386 147084 185686
<< nwell >>
rect 21084 185436 147184 185786
rect 21084 30636 21434 185436
rect 146834 30636 147184 185436
rect 21084 30286 147184 30636
<< nsubdiff >>
rect 21184 185686 21284 185711
rect 146984 185686 147084 185711
rect 21159 185586 21284 185686
rect 146984 185586 147109 185686
rect 21184 185536 21284 185586
rect 21184 30486 21284 30536
rect 146984 185536 147084 185586
rect 146984 30486 147084 30536
rect 21159 30386 21284 30486
rect 146984 30386 147109 30486
rect 21184 30361 21284 30386
rect 146984 30361 147084 30386
<< nsubdiffcont >>
rect 21284 185586 146984 185686
rect 21184 30536 21284 185536
rect 146984 30536 147084 185536
rect 21284 30386 146984 30486
<< locali >>
rect 21134 185686 147134 185736
rect 21134 185586 21284 185686
rect 146984 185586 147134 185686
rect 21134 185536 147134 185586
rect 21134 30536 21184 185536
rect 21284 30536 21334 185536
rect 146934 30536 146984 185536
rect 147084 30536 147134 185536
rect 21134 30486 147134 30536
rect 21134 30386 21284 30486
rect 146984 30386 147134 30486
rect 21134 30336 147134 30386
<< metal2 >>
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect -800 680242 1700 685242
rect 582300 677984 584800 682984
rect -800 643842 1660 648642
rect 582340 639784 584800 644584
rect -800 633842 1660 638642
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use sonos_array_50x50x64  sonos_array_50x50x64_0
timestamp 1685137779
transform 1 0 21694 0 1 30912
box -80 -96 125116 154280
use sonos_array_labeled  sonos_array_labeled_0
array 0 19 14496 0 19 15060
timestamp 1685135448
transform 1 0 179200 0 1 38600
box 0 0 4496 5060
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
