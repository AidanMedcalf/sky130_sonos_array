magic
tech sky130A
timestamp 1686079789
<< error_p >>
rect -72 109 72 174
rect 72 -126 228 109
<< dnwell >>
rect -72 -126 72 109
<< npd >>
rect -45 21 45 51
<< nsonos >>
rect -45 -65 45 -21
<< ndiff >>
rect -45 93 45 101
rect -45 59 -17 93
rect 17 59 45 93
rect -45 51 45 59
rect -45 -21 45 21
rect -45 -80 45 -65
rect -45 -114 -17 -80
rect 17 -114 45 -80
rect -45 -122 45 -114
<< ndiffc >>
rect -17 59 17 93
rect -17 -114 17 -80
<< poly >>
rect -72 21 -45 51
rect 45 21 72 51
rect -72 -65 -45 -21
rect 45 -65 72 -21
<< locali >>
rect -22 93 88 109
rect -22 59 -17 93
rect 17 59 53 93
rect 87 59 88 93
rect -22 43 88 59
rect -72 -30 72 4
rect -33 -80 33 -72
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -122 33 -114
<< viali >>
rect 53 59 87 93
rect -17 -114 17 -80
<< metal1 >>
rect -18 -74 18 101
rect 52 99 88 105
rect 47 93 93 99
rect 47 59 53 93
rect 87 59 93 93
rect 47 53 93 59
rect -23 -80 23 -74
rect -23 -114 -17 -80
rect 17 -114 23 -80
rect -23 -120 23 -114
rect -18 -126 18 -120
rect 52 -122 88 53
<< properties >>
string FIXED_BBOX -72 -126 93 109
<< end >>
