magic
tech sky130A
timestamp 1686033482
<< error_s >>
rect -80 1387 1250 1530
rect -80 1381 63 1387
rect 1107 1381 1250 1387
rect -80 1337 117 1381
rect 171 1337 261 1381
rect 315 1337 405 1381
rect 459 1337 549 1381
rect 603 1337 693 1381
rect 747 1337 837 1381
rect 891 1337 981 1381
rect 1035 1337 1250 1381
rect -80 1143 63 1337
rect 1107 1143 1250 1337
rect -80 1099 117 1143
rect 171 1099 261 1143
rect 315 1099 405 1143
rect 459 1099 549 1143
rect 603 1099 693 1143
rect 747 1099 837 1143
rect 891 1099 981 1143
rect 1035 1099 1250 1143
rect -80 1035 63 1099
rect 1107 1035 1250 1099
rect -80 991 117 1035
rect 171 991 261 1035
rect 315 991 405 1035
rect 459 991 549 1035
rect 603 991 693 1035
rect 747 991 837 1035
rect 891 991 981 1035
rect 1035 991 1250 1035
rect -80 797 63 991
rect 1107 797 1250 991
rect -80 753 117 797
rect 171 753 261 797
rect 315 753 405 797
rect 459 753 549 797
rect 603 753 693 797
rect 747 753 837 797
rect 891 753 981 797
rect 1035 753 1250 797
rect -80 689 63 753
rect 1107 689 1250 753
rect -80 645 117 689
rect 171 645 261 689
rect 315 645 405 689
rect 459 645 549 689
rect 603 645 693 689
rect 747 645 837 689
rect 891 645 981 689
rect 1035 645 1250 689
rect -80 451 63 645
rect 1107 451 1250 645
rect -80 407 117 451
rect 171 407 261 451
rect 315 407 405 451
rect 459 407 549 451
rect 603 407 693 451
rect 747 407 837 451
rect 891 407 981 451
rect 1035 407 1250 451
rect -80 343 63 407
rect 1107 343 1250 407
rect -80 299 117 343
rect 171 299 261 343
rect 315 299 405 343
rect 459 299 549 343
rect 603 299 693 343
rect 747 299 837 343
rect 891 299 981 343
rect 1035 299 1250 343
rect -80 105 63 299
rect 1107 105 1250 299
rect -80 61 117 105
rect 171 61 261 105
rect 315 61 405 105
rect 459 61 549 105
rect 603 61 693 105
rect 747 61 837 105
rect 891 61 981 105
rect 1035 61 1250 105
rect -80 55 63 61
rect 1107 55 1250 61
rect -80 -88 1250 55
<< dnwell >>
rect -40 -48 1210 1490
<< psubdiff >>
rect -40 1486 1210 1490
rect -40 1469 0 1486
rect 1173 1469 1210 1486
rect -40 1465 1210 1469
rect -40 1438 -15 1465
rect -40 4 -36 1438
rect -19 4 -15 1438
rect 1185 1438 1210 1465
rect -40 -23 -15 4
rect 1185 4 1189 1438
rect 1206 4 1210 1438
rect 1185 -23 1210 4
rect -40 -27 1210 -23
rect -40 -44 0 -27
rect 1173 -44 1210 -27
rect -40 -48 1210 -44
<< psubdiffcont >>
rect 0 1469 1173 1486
rect -36 4 -19 1438
rect 1189 4 1206 1438
rect 0 -44 1173 -27
<< poly >>
rect 1140 1370 1173 1381
rect 1140 1346 1144 1370
rect 1161 1346 1173 1370
rect 1140 1292 1173 1346
rect 1140 1268 1144 1292
rect 1161 1268 1173 1292
rect 1140 1212 1173 1268
rect 1140 1188 1144 1212
rect 1161 1188 1173 1212
rect 1140 1132 1173 1188
rect 1140 1108 1144 1132
rect 1161 1108 1173 1132
rect 1140 1025 1173 1108
rect 1140 1001 1144 1025
rect 1161 1001 1173 1025
rect 1140 946 1173 1001
rect 1140 922 1144 946
rect 1161 922 1173 946
rect 1140 866 1173 922
rect 1140 842 1144 866
rect 1161 842 1173 866
rect 1140 787 1173 842
rect 1140 763 1144 787
rect 1161 763 1173 787
rect 1140 679 1173 763
rect 1140 655 1144 679
rect 1161 655 1173 679
rect 1140 600 1173 655
rect 1140 576 1144 600
rect 1161 576 1173 600
rect 1140 520 1173 576
rect 1140 496 1144 520
rect 1161 496 1173 520
rect 1140 440 1173 496
rect 1140 416 1144 440
rect 1161 416 1173 440
rect 1140 333 1173 416
rect 1140 309 1144 333
rect 1161 309 1173 333
rect 1140 254 1173 309
rect 1140 230 1144 254
rect 1161 230 1173 254
rect 1140 174 1173 230
rect 1140 150 1144 174
rect 1161 150 1173 174
rect 1140 97 1173 150
rect 1140 73 1144 97
rect 1161 73 1173 97
rect 1140 61 1173 73
<< polycont >>
rect 1144 1346 1161 1370
rect 1144 1268 1161 1292
rect 1144 1188 1161 1212
rect 1144 1108 1161 1132
rect 1144 1001 1161 1025
rect 1144 922 1161 946
rect 1144 842 1161 866
rect 1144 763 1161 787
rect 1144 655 1161 679
rect 1144 576 1161 600
rect 1144 496 1161 520
rect 1144 416 1161 440
rect 1144 309 1161 333
rect 1144 230 1161 254
rect 1144 150 1161 174
rect 1144 73 1161 97
<< locali >>
rect -36 1469 0 1486
rect 1173 1469 1206 1486
rect -36 1438 -19 1469
rect 39 1438 1113 1469
rect 1189 1438 1206 1469
rect 1136 1370 1189 1381
rect 1136 1346 1144 1370
rect 1161 1346 1189 1370
rect -19 1312 0 1346
rect 1136 1292 1189 1346
rect 1136 1268 1144 1292
rect 1161 1268 1189 1292
rect 1136 1212 1189 1268
rect 1136 1188 1144 1212
rect 1161 1188 1189 1212
rect -19 1134 0 1168
rect 1136 1132 1189 1188
rect 1136 1108 1144 1132
rect 1161 1108 1189 1132
rect 1136 1025 1189 1108
rect 1136 1001 1144 1025
rect 1161 1001 1189 1025
rect -19 966 0 1000
rect 1136 946 1189 1001
rect 1136 922 1144 946
rect 1161 922 1189 946
rect 1136 866 1189 922
rect 1136 842 1144 866
rect 1161 842 1189 866
rect -19 788 0 822
rect 1136 787 1189 842
rect 1136 763 1144 787
rect 1161 763 1189 787
rect 1136 679 1189 763
rect 1136 655 1144 679
rect 1161 655 1189 679
rect -19 620 0 654
rect 1136 600 1189 655
rect 1136 576 1144 600
rect 1161 576 1189 600
rect 1136 520 1189 576
rect 1136 496 1144 520
rect 1161 496 1189 520
rect -19 442 0 476
rect 1136 440 1189 496
rect 1136 416 1144 440
rect 1161 416 1189 440
rect 1136 333 1189 416
rect 1136 309 1144 333
rect 1161 309 1189 333
rect -19 274 0 308
rect 1136 254 1189 309
rect 1136 230 1144 254
rect 1161 230 1189 254
rect 1136 174 1189 230
rect 1136 150 1144 174
rect 1161 150 1189 174
rect -19 96 0 130
rect 1136 97 1189 150
rect 1136 73 1144 97
rect 1161 73 1189 97
rect 1136 61 1189 73
rect -36 -27 -19 4
rect 39 -27 1113 4
rect 1189 -27 1206 4
rect -36 -44 0 -27
rect 1173 -44 1206 -27
<< metal1 >>
rect 95 1390 1152 1436
rect 92 6 1155 52
use sonos_cell_mirrored  sonos_cell_mirrored_0
array 0 7 144 0 3 346
timestamp 1686033482
transform 1 0 -80 0 1 -80
box 40 40 380 524
<< end >>
