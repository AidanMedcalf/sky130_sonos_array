magic
tech sky130A
timestamp 1663450679
<< error_p >>
rect 0 566 165 699
rect -40 526 205 566
rect -40 399 300 526
rect -40 359 205 399
<< dnwell >>
rect 0 399 165 526
<< psubdiff >>
rect 0 514 165 526
rect 0 489 24 514
rect 141 489 165 514
rect 0 477 165 489
<< psubdiffcont >>
rect 24 489 141 514
<< metal1 >>
rect 0 412 165 458
rect 54 404 90 412
rect 124 400 160 412
<< end >>
