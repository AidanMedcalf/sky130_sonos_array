magic
tech sky130A
timestamp 1686033289
<< error_p >>
rect -502 -152 40 -130
rect -530 -170 40 -152
rect -512 -188 -467 -170
rect -249 -465 40 -170
rect 0 -683 40 -465
rect -18 -718 40 -683
rect -18 -728 18 -718
rect 0 -746 18 -728
<< dnwell >>
rect -462 -678 0 -170
<< nwell >>
rect -548 -465 -249 -170
rect -548 -764 0 -465
<< srampvar >>
rect -111 -276 -36 -246
<< psubdiff >>
rect -111 -246 -36 -170
rect -111 -362 -36 -276
rect -111 -438 0 -362
<< nsubdiff >>
rect -512 -212 -467 -170
rect -512 -524 -507 -212
rect -473 -524 -467 -212
rect -512 -683 -467 -524
rect -512 -689 0 -683
rect -512 -723 -309 -689
rect -18 -723 0 -689
rect -512 -728 0 -723
<< nsubdiffcont >>
rect -507 -524 -473 -212
rect -309 -723 -18 -689
<< poly >>
rect -25 -246 5 -216
rect -203 -263 -111 -246
rect -203 -297 -193 -263
rect -159 -276 -111 -263
rect -36 -276 5 -246
rect -159 -297 -149 -276
rect -203 -313 -149 -297
<< polycont >>
rect -193 -297 -159 -263
<< locali >>
rect -507 -212 -473 -170
rect -91 -263 -57 -223
rect -209 -297 -193 -263
rect -159 -278 -57 -263
rect -159 -297 -91 -278
rect -91 -380 -57 -312
rect -106 -414 -91 -380
rect -57 -414 0 -380
rect -91 -430 -57 -414
rect -507 -689 -473 -524
rect -507 -723 -309 -689
rect -18 -723 0 -689
<< viali >>
rect -91 -312 -57 -278
rect -91 -414 -57 -380
<< metal1 >>
rect -111 -278 -50 -170
rect -111 -312 -91 -278
rect -57 -312 -50 -278
rect -111 -380 -50 -312
rect -111 -414 -91 -380
rect -57 -414 -50 -380
rect -111 -438 -50 -414
<< end >>
