magic
tech sky130A
timestamp 1663450679
<< error_p >>
rect -152 404 73 444
rect -152 0 188 404
rect -152 -40 73 0
<< dnwell >>
rect -112 0 33 404
<< psubdiff >>
rect -112 346 -63 404
rect -112 58 -100 346
rect -75 58 -63 346
rect -112 0 -63 58
<< psubdiffcont >>
rect -100 58 -75 346
<< poly >>
rect -44 343 0 346
rect -44 338 33 343
rect -44 304 -39 338
rect -5 304 33 338
rect -44 299 33 304
rect -44 257 0 299
rect -44 252 33 257
rect -44 232 -39 252
rect -5 232 33 252
rect -44 227 33 232
rect -44 177 0 227
rect -44 172 33 177
rect -44 152 -39 172
rect -5 152 33 172
rect -44 147 33 152
rect -44 104 0 147
rect -44 100 33 104
rect -44 66 -39 100
rect -5 66 33 100
rect -44 61 33 66
rect -44 58 0 61
<< polycont >>
rect -39 304 -5 338
rect -39 232 -5 252
rect -39 152 -5 172
rect -39 66 -5 100
<< locali >>
rect -44 338 0 404
rect -44 304 -39 338
rect -5 304 0 338
rect -44 252 0 304
rect -44 232 -39 252
rect -5 232 0 252
rect -44 172 0 232
rect -44 152 -39 172
rect -5 152 0 172
rect -44 100 0 152
rect -44 66 -39 100
rect -5 66 0 100
rect -44 0 0 66
<< end >>
