magic
tech sky130A
timestamp 1685642023
<< dnwell >>
rect -2800 1800 2800 3800
<< nwell >>
rect -2860 3690 2860 3860
rect -2860 1910 -2690 3690
rect 2690 1910 2860 3690
rect -2860 1740 2860 1910
<< pwell >>
rect -3050 3860 3050 4050
rect -3050 1740 -2860 3860
rect 2860 1740 3050 3860
rect -3050 1550 3050 1740
<< mvpsubdiff >>
rect -3000 3910 -2800 4000
rect 2660 3910 3000 4000
rect -3000 3810 -2910 3910
rect -3000 1690 -2910 1800
rect 2910 3810 3000 3910
rect 2910 1690 3000 1800
rect -3000 1600 -2800 1690
rect 2660 1600 3000 1690
<< mvnsubdiff >>
rect -2820 3730 -2650 3820
rect 2650 3730 2820 3820
rect -2820 3650 -2730 3730
rect -2820 1870 -2730 1950
rect 2730 3650 2820 3730
rect 2730 1870 2820 1950
rect -2820 1780 -2650 1870
rect 2650 1780 2820 1870
<< mvpsubdiffcont >>
rect -2800 3910 2660 4000
rect -3000 1800 -2910 3810
rect 2910 1800 3000 3810
rect -2800 1600 2660 1690
<< mvnsubdiffcont >>
rect -2650 3730 2650 3820
rect -2820 1950 -2730 3650
rect 2730 1950 2820 3650
rect -2650 1780 2650 1870
<< locali >>
rect -3000 3910 -2800 4000
rect 2660 3910 3000 4000
rect -3000 3810 -2910 3910
rect -3000 1690 -2910 1800
rect -2820 3730 -2650 3820
rect 2650 3730 2820 3820
rect -2820 3650 -2730 3730
rect -2820 1870 -2730 1950
rect 2730 3650 2820 3730
rect 2730 1870 2820 1950
rect -2820 1780 -2650 1870
rect 2650 1780 2820 1870
rect 2910 3810 3000 3910
rect 2910 1690 3000 1800
rect -3000 1600 -2800 1690
rect 2660 1600 3000 1690
<< metal1 >>
rect -3000 3910 3000 4000
rect -3000 1690 -2910 3910
rect -2820 3730 2820 3820
rect -2820 1870 -2730 3730
rect 2730 1870 2820 3730
rect -2820 1780 2820 1870
rect 2910 1690 3000 3910
rect -3000 1600 3000 1690
use sky130_ef_io__esd_pdiode_11v0_array  sky130_ef_io__esd_pdiode_11v0_array_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1685637275
transform 0 1 -6 -1 0 2783
box -783 -2594 783 2594
use tp_pad_m5  tp_pad_m5_0
timestamp 1685412872
transform 1 0 0 0 1 2000
box -2000 -2000 2000 2000
<< end >>
