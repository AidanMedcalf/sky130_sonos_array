* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_5p73_JY438B a_n573_50# a_n573_n482# w_n802_n711#
+ VSUBS
X0 a_n573_50# a_n573_n482# VSUBS sky130_fd_pr__res_xhigh_po w=5.73 l=0.5
.ends

.subckt sky130_fd_bs_flash__special_sonosfet_star w_n436_n442# a_n33_36# dw_n436_n442#
+ a_22_n76# a_n84_n76#
X0 a_22_n76# a_n33_36# a_n84_n76# w_n436_n442# sky130_fd_bs_flash__special_sonosfet_star ad=0.14 pd=1.52 as=0.14 ps=1.52 w=0.45 l=0.22
.ends

.subckt sonos_1t_iso G D VNB S B
Xsky130_fd_bs_flash__special_sonosfet_star_0 B G VNB D S sky130_fd_bs_flash__special_sonosfet_star
.ends

.subckt sonos_endcap_tb dw_n408_n1786# m1_n300_n1886# w_n120_n1786# w_n408_n1360#
+ a_n408_n922# a_n354_n1046#
X0 a_n354_n1046# a_n408_n922# a_n354_n1046# w_n408_n1360# sky130_fd_pr__nfet_01v8 ad=1.01 pd=5.84 as=0.45 ps=2.8 w=0.9 l=0.3
.ends

.subckt sonos_cell w_n144_n252# a_n144_n130# dw_n144_n252# a_n90_n244# a_n90_102#
+ li_n144_n60# a_n144_42#
X0 a_n90_102# a_n144_42# a_n90_n42# w_n144_n252# sky130_fd_pr__special_nfet_latch ad=0.45 pd=2.8 as=0.189 ps=1.32 w=0.9 l=0.3
X1 a_n90_n42# a_n144_n130# a_n90_n244# w_n144_n252# sky130_fd_bs_flash__special_sonosfet_star ad=0.189 pd=1.32 as=0.513 ps=2.94 w=0.9 l=0.44
.ends

.subckt sonos_array_orig sonos_endcap_lr_1[3]/a_n616_n202# sonos_endcap_lr_1[0]/a_n454_n406#
+ sonos_cell_2[2|7]/li_n144_n60# sonos_endcap_lr_2[1]/a_n616_n202# sonos_endcap_lr_2[0]/a_n616_28#
+ sonos_endcap_lr_1[3]/a_n454_n406# sonos_endcap_lr_2[1]/a_n616_28# sonos_endcap_lr_2[1]/a_n454_n406#
+ sonos_endcap_lr_2[2]/a_n616_28# sonos_endcap_lr_2[3]/a_n616_28# sonos_endcap_lr_1[1]/a_n616_n202#
+ sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|4]/a_n90_102# sonos_endcap_lr_1[1]/a_n454_n406#
+ sonos_cell_1[3|7]/li_n144_n60# sonos_cell_2[3|1]/a_n90_n244# sonos_endcap_lr_2[2]/a_n616_n202#
+ sonos_cell_2[3|6]/a_n90_n244# sonos_endcap_lr_2[2]/a_n454_n406# sonos_cell_2[3|1]/a_n90_102#
+ sonos_cell_1[2|7]/li_n144_n60# sonos_cell_2[3|0]/a_n90_n244# sonos_endcap_lr_1[2]/a_n616_n202#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[3|3]/a_n90_n244#
+ dw_0_n64# sonos_cell_2[3|5]/a_n90_n244# sonos_endcap_lr_2[0]/a_n616_n202# sonos_cell_2[3|3]/a_n90_102#
+ w_n498_n930# sonos_endcap_lr_1[2]/a_n454_n406# sonos_endcap_lr_1[0]/a_n616_28# sonos_cell_2[3|7]/a_n90_102#
+ sonos_endcap_lr_1[1]/a_n616_28# sonos_cell_1[1|7]/li_n144_n60# sonos_endcap_lr_2[3]/a_n616_n202#
+ sonos_endcap_lr_1[2]/a_n616_28# sonos_cell_2[3|4]/a_n90_n244# sonos_endcap_lr_2[0]/a_n454_n406#
+ sonos_endcap_lr_1[3]/a_n616_28# sonos_cell_2[3|2]/a_n90_102# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_endcap_lr_1[0]/a_n616_n202# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_1[0|7]/li_n144_n60# sonos_cell_2[3|0]/a_n90_102#
+ sonos_endcap_lr_2[3]/a_n454_n406#
Xsonos_endcap_tb_1[0] dw_0_n64# sonos_cell_2[3|0]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|0]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[1] dw_0_n64# sonos_cell_2[3|1]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|1]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[2] dw_0_n64# sonos_cell_2[3|2]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|2]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[3] dw_0_n64# sonos_cell_2[3|3]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|3]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[4] dw_0_n64# sonos_cell_2[3|4]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|4]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[5] dw_0_n64# sonos_cell_2[3|5]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|5]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[6] dw_0_n64# sonos_cell_2[3|6]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|6]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[7] dw_0_n64# sonos_cell_2[3|7]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|7]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[0] dw_0_n64# sonos_cell_2[3|0]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|0]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[1] dw_0_n64# sonos_cell_2[3|1]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|1]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[2] dw_0_n64# sonos_cell_2[3|2]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|2]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[3] dw_0_n64# sonos_cell_2[3|3]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|3]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[4] dw_0_n64# sonos_cell_2[3|4]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|4]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[5] dw_0_n64# sonos_cell_2[3|5]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|5]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[6] dw_0_n64# sonos_cell_2[3|6]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|6]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[7] dw_0_n64# sonos_cell_2[3|7]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|7]/a_n90_102# sonos_endcap_tb
Xsonos_cell_1[0|0] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244# sonos_cell_2[3|0]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|0] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|0] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|0] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|1] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244# sonos_cell_2[3|1]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|1] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|1] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|1] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|2] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244# sonos_cell_2[3|2]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|2] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|2] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|2] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|3] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244# sonos_cell_2[3|3]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|3] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|3] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|3] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|4] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244# sonos_cell_2[3|4]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|4] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|4] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|4] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|5] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244# sonos_cell_2[3|5]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|5] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|5] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|5] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|6] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244# sonos_cell_2[3|6]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|6] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|6] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|6] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|7] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244# sonos_cell_2[3|7]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|7] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|7] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|7] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|0] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|0] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|0] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|0] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|1] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|1] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|1] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|1] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|2] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|2] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|2] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|2] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|3] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|3] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|3] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|3] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|4] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|4] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|4] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|4] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|5] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|5] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|5] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|5] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|6] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|6] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|6] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|6] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|7] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|7] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|7] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|7] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
.ends

.subckt sonos_array_labeled WL2 WL1 WL0 PT7 PT6 PT5 PT4 PT3 PT2 PT1 PT0 VPB WLS7 WLS6
+ BL2 WLS5 BL1 WLS4 BL0 WLS3 WLS2 WLS1 WLS0 VNB SRC2 SRC1 SRC0
Xsonos_array_orig_0 WLS1 WL7 PT3 WLS2 WLS1 WL1 WLS3 WL2 WLS5 WLS7 WLS5 PT1 SRC4 WL5
+ PT0 BL1 WLS4 BL6 WL4 SRC1 PT2 BL0 WLS3 SRC5 PT7 BL3 VNB BL5 WLS0 SRC3 VPB WL3 WLS6
+ SRC7 WLS4 PT4 WLS6 WLS2 BL4 WL0 WLS0 SRC2 BL2 WLS7 PT5 BL7 SRC6 PT6 SRC0 WL6 sonos_array_orig
.ends

.subckt sonos_cell_mirrored sonos_cell_0/a_n144_n130# sonos_cell_0/a_n144_42# w_160_160#
+ sonos_cell_1/a_n144_42# sonos_cell_0/li_n144_n60# sonos_cell_1/a_n90_102# sonos_cell_1/dw_n144_n252#
+ sonos_cell_1/a_n144_n130# sonos_cell_1/a_n90_n244# sonos_cell_1/li_n144_n60#
Xsonos_cell_0 w_160_160# sonos_cell_0/a_n144_n130# sonos_cell_1/dw_n144_n252# sonos_cell_1/a_n90_n244#
+ sonos_cell_1/a_n90_102# sonos_cell_0/li_n144_n60# sonos_cell_0/a_n144_42# sonos_cell
Xsonos_cell_1 w_160_160# sonos_cell_1/a_n144_n130# sonos_cell_1/dw_n144_n252# sonos_cell_1/a_n90_n244#
+ sonos_cell_1/a_n90_102# sonos_cell_1/li_n144_n60# sonos_cell_1/a_n144_42# sonos_cell
.ends

.subckt sonos_8x8 w_n80_n96# dw_n80_n96#
Xsonos_cell_mirrored_0[0|0] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|0] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|0] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|0] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|1] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|1] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|1] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|1] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|2] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|2] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|2] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|2] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|3] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|3] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|3] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|3] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|4] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|4] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|4] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|4] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|5] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|5] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|5] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|5] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|6] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|6] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|6] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|6] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|7] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|7] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|7] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|7] w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
.ends

.subckt sonos_array_1x1x64 w_n80_n96# dw_n80_n96#
Xsonos_8x8_0 w_n80_n96# dw_n80_n96# sonos_8x8
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_8 m1_379680_149580# sonos_1t_iso_7/B li_379366_150034#
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_9 m1_367680_149580# D li_367366_150034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_1t_iso_11 G D sonos_1t_iso_11/VNB S sonos_1t_iso_11/B sonos_1t_iso
Xsonos_1t_iso_10 G D sonos_1t_iso_10/VNB S sonos_1t_iso_10/B sonos_1t_iso
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_20 m1_427680_149580# G li_427366_150034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_1t_iso_12 G D sonos_1t_iso_12/VNB S sonos_1t_iso_12/B sonos_1t_iso
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_21 m1_415680_149580# S sonos_1t_iso_15/VNB
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_10 m1_355680_149580# G li_355366_150034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_1t_iso_13 G D sonos_1t_iso_13/VNB S sonos_1t_iso_13/B sonos_1t_iso
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_22 m1_451680_165580# sonos_1t_iso_14/B li_451366_166034#
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_1t_iso_14 G D sonos_1t_iso_14/VNB S sonos_1t_iso_14/B sonos_1t_iso
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_23 m1_451680_149580# sonos_1t_iso_15/B li_451366_150034#
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_12 m1_415680_133580# S sonos_1t_iso_13/VNB
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_11 m1_343680_149580# S sonos_1t_iso_7/VNB
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_13 m1_427680_133580# G li_427366_134034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_1t_iso_15 G D sonos_1t_iso_15/VNB S sonos_1t_iso_15/B sonos_1t_iso
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_14 m1_439680_133580# D li_439366_134034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_15 m1_451680_133580# sonos_1t_iso_13/B li_451366_134034#
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_16 m1_415680_165580# S sonos_1t_iso_14/VNB
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_17 m1_427680_165580# G li_427366_166034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_18 m1_439680_165580# D li_439366_166034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_19 m1_439680_149580# D li_439366_150034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_1t_iso_0 sonos_1t_iso_0/G sonos_1t_iso_0/D sonos_1t_iso_0/VNB sonos_1t_iso_0/S
+ sonos_1t_iso_0/B sonos_1t_iso
Xsonos_1t_iso_1 G D sonos_1t_iso_1/VNB S sonos_1t_iso_1/B sonos_1t_iso
Xsonos_1t_iso_2 G D sonos_1t_iso_2/VNB S sonos_1t_iso_2/B sonos_1t_iso
Xsonos_1t_iso_3 G D sonos_1t_iso_3/VNB S sonos_1t_iso_3/B sonos_1t_iso
Xsonos_1t_iso_4 G D sonos_1t_iso_4/VNB S sonos_1t_iso_4/B sonos_1t_iso
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_0 m1_367680_165580# D li_367366_166034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_1t_iso_5 G D sonos_1t_iso_5/VNB S sonos_1t_iso_5/B sonos_1t_iso
Xsonos_1t_iso_6 G D sonos_1t_iso_6/VNB S sonos_1t_iso_6/B sonos_1t_iso
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_2 m1_355680_133580# G li_355366_134034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_1 m1_367680_133580# D li_367366_134034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_1t_iso_7 G D sonos_1t_iso_7/VNB S sonos_1t_iso_7/B sonos_1t_iso
Xsonos_array_labeled_0 sonos_array_labeled_0/WL2 sonos_array_labeled_0/WL1 sonos_array_labeled_0/WL0
+ sonos_array_labeled_0/PT7 sonos_array_labeled_0/PT6 sonos_array_labeled_0/PT5 sonos_array_labeled_0/PT4
+ sonos_array_labeled_0/PT3 sonos_array_labeled_0/PT2 sonos_array_labeled_0/PT1 sonos_array_labeled_0/PT0
+ sonos_array_labeled_0/VPB sonos_array_labeled_0/PT7 sonos_array_labeled_0/PT6 sonos_array_labeled_0/BL2
+ sonos_array_labeled_0/PT5 sonos_array_labeled_0/BL1 sonos_array_labeled_0/PT4 sonos_array_labeled_0/BL0
+ sonos_array_labeled_0/PT3 sonos_array_labeled_0/PT2 sonos_array_labeled_0/PT1 sonos_array_labeled_0/PT0
+ sonos_array_labeled_0/VNB sonos_array_labeled_0/SRC2 sonos_array_labeled_0/SRC1
+ sonos_array_labeled_0/SRC0 sonos_array_labeled
Xsonos_array_1x1x64_0[0|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|0] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|1] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|2] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|3] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|4] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|5] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|6] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|7] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|8] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|9] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|10] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|11] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|12] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|13] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|14] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|15] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|16] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|17] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|18] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|19] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|20] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|21] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|22] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|23] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[0|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[1|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[2|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[3|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[4|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[5|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[6|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[7|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[8|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[9|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[10|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[11|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[12|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[13|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[14|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[15|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[16|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[17|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[18|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[19|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[20|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[21|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[22|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[23|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[24|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[25|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[26|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[27|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[28|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsonos_array_1x1x64_0[29|24] w_229206_435606# dw_229000_435400# sonos_array_1x1x64
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_3 m1_379680_165580# sonos_1t_iso_6/B li_379366_166034#
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_array_labeled_1 sonos_array_labeled_1/WL2 sonos_array_labeled_1/WL1 sonos_array_labeled_1/WL0
+ sonos_array_labeled_1/PT7 sonos_array_labeled_1/PT6 sonos_array_labeled_1/PT5 sonos_array_labeled_1/PT4
+ sonos_array_labeled_1/PT3 sonos_array_labeled_1/PT2 sonos_array_labeled_1/PT1 sonos_array_labeled_1/PT0
+ sonos_array_labeled_1/VPB sonos_array_labeled_1/PT7 sonos_array_labeled_1/PT6 sonos_array_labeled_1/BL2
+ sonos_array_labeled_1/PT5 sonos_array_labeled_1/BL1 sonos_array_labeled_1/PT4 sonos_array_labeled_1/BL0
+ sonos_array_labeled_1/PT3 sonos_array_labeled_1/PT2 sonos_array_labeled_1/PT1 sonos_array_labeled_1/PT0
+ sonos_array_labeled_1/VNB sonos_array_labeled_1/SRC2 sonos_array_labeled_1/SRC1
+ sonos_array_labeled_1/SRC0 sonos_array_labeled
Xsonos_1t_iso_8 sonos_1t_iso_8/G sonos_1t_iso_8/D sonos_1t_iso_8/VNB sonos_1t_iso_8/S
+ sonos_1t_iso_8/B sonos_1t_iso
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_4 m1_343680_133580# S sonos_1t_iso_1/VNB vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_array_labeled_2 sonos_array_labeled_2/WL2 sonos_array_labeled_2/WL1 sonos_array_labeled_2/WL0
+ sonos_array_labeled_2/PT7 sonos_array_labeled_2/PT6 sonos_array_labeled_2/PT5 sonos_array_labeled_2/PT4
+ sonos_array_labeled_2/PT3 sonos_array_labeled_2/PT2 sonos_array_labeled_2/PT1 sonos_array_labeled_2/PT0
+ sonos_array_labeled_2/VPB sonos_array_labeled_2/PT7 sonos_array_labeled_2/PT6 sonos_array_labeled_2/BL2
+ sonos_array_labeled_2/PT5 sonos_array_labeled_2/BL1 sonos_array_labeled_2/PT4 sonos_array_labeled_2/BL0
+ sonos_array_labeled_2/PT3 sonos_array_labeled_2/PT2 sonos_array_labeled_2/PT1 sonos_array_labeled_2/PT0
+ sonos_array_labeled_2/VNB sonos_array_labeled_2/SRC2 sonos_array_labeled_2/SRC1
+ sonos_array_labeled_2/SRC0 sonos_array_labeled
Xsonos_1t_iso_9 G D sonos_1t_iso_9/VNB S sonos_1t_iso_9/B sonos_1t_iso
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_5 m1_355680_165580# G li_355366_166034# vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_array_labeled_3 sonos_array_labeled_3/WL2 sonos_array_labeled_3/WL1 sonos_array_labeled_3/WL0
+ sonos_array_labeled_3/PT7 sonos_array_labeled_3/PT6 sonos_array_labeled_3/PT5 sonos_array_labeled_3/PT4
+ sonos_array_labeled_3/PT3 sonos_array_labeled_3/PT2 sonos_array_labeled_3/PT1 sonos_array_labeled_3/PT0
+ sonos_array_labeled_3/VPB sonos_array_labeled_3/PT7 sonos_array_labeled_3/PT6 sonos_array_labeled_3/BL2
+ sonos_array_labeled_3/PT5 sonos_array_labeled_3/BL1 sonos_array_labeled_3/PT4 sonos_array_labeled_3/BL0
+ sonos_array_labeled_3/PT3 sonos_array_labeled_3/PT2 sonos_array_labeled_3/PT1 sonos_array_labeled_3/PT0
+ sonos_array_labeled_3/VNB sonos_array_labeled_3/SRC2 sonos_array_labeled_3/SRC1
+ sonos_array_labeled_3/SRC0 sonos_array_labeled
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_6 m1_343680_165580# S sonos_1t_iso_6/VNB vssa1
+ sky130_fd_pr__res_xhigh_po_5p73_JY438B
Xsonos_array_labeled_4 sonos_array_labeled_4/WL2 sonos_array_labeled_4/WL1 sonos_array_labeled_4/WL0
+ sonos_array_labeled_4/PT7 sonos_array_labeled_4/PT6 sonos_array_labeled_4/PT5 sonos_array_labeled_4/PT4
+ sonos_array_labeled_4/PT3 sonos_array_labeled_4/PT2 sonos_array_labeled_4/PT1 sonos_array_labeled_4/PT0
+ sonos_array_labeled_4/VPB sonos_array_labeled_4/PT7 sonos_array_labeled_4/PT6 sonos_array_labeled_4/BL2
+ sonos_array_labeled_4/PT5 sonos_array_labeled_4/BL1 sonos_array_labeled_4/PT4 sonos_array_labeled_4/BL0
+ sonos_array_labeled_4/PT3 sonos_array_labeled_4/PT2 sonos_array_labeled_4/PT1 sonos_array_labeled_4/PT0
+ sonos_array_labeled_4/VNB sonos_array_labeled_4/SRC2 sonos_array_labeled_4/SRC1
+ sonos_array_labeled_4/SRC0 sonos_array_labeled
Xsky130_fd_pr__res_xhigh_po_5p73_JY438B_7 m1_379680_133580# sonos_1t_iso_1/B li_379366_134034#
+ vssa1 sky130_fd_pr__res_xhigh_po_5p73_JY438B
.ends

