magic
tech sky130A
timestamp 1686079789
<< dnwell >>
rect 0 -32 1 177
<< nwell >>
rect 1569 -633 1608 1635
<< poly >>
rect 0 100 1 130
rect 0 14 1 58
use sonos_array_corner  sonos_array_corner_1
timestamp 1686079789
transform 1 0 0 0 1 0
box -548 -764 18 -152
use sonos_array_corner  sonos_array_corner_2
timestamp 1686079789
transform 1 0 0 0 -1 1002
box -548 -764 18 -152
use sonos_array_corner  sonos_array_corner_3
timestamp 1686079789
transform -1 0 1152 0 1 0
box -548 -764 18 -152
use sonos_array_corner  sonos_array_corner_4
timestamp 1686079789
transform -1 0 1152 0 -1 1002
box -548 -764 18 -152
use sonos_cell  sonos_cell_1
array 0 7 144 0 3 346
timestamp 1686079789
transform 1 0 72 0 1 79
box -72 -126 228 174
use sonos_cell  sonos_cell_2
array 0 7 144 0 3 -346
timestamp 1686079789
transform 1 0 72 0 -1 -115
box -72 -126 228 174
use sonos_endcap_lr  sonos_endcap_lr_1
array 0 0 417 0 3 346
timestamp 1686079789
transform 1 0 0 0 1 0
box -548 -230 0 152
use sonos_endcap_lr  sonos_endcap_lr_2
array 0 0 417 0 3 346
timestamp 1686079789
transform -1 0 1152 0 -1 1002
box -548 -230 0 152
use sonos_endcap_tb  sonos_endcap_tb_1
array 0 7 144 0 0 154
timestamp 1686079789
transform 1 0 204 0 1 215
box -222 -979 96 -373
use sonos_endcap_tb  sonos_endcap_tb_2
array 0 7 144 0 0 -154
timestamp 1686079789
transform 1 0 204 0 -1 787
box -222 -979 96 -373
<< end >>
