* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sonos_cell w_n144_n252# a_n144_n130# dw_n144_n252# a_n90_n244# a_n90_102#
+ li_n144_n60# a_n144_42#
X0 a_n90_102# a_n144_42# a_n90_n42# w_n144_n252# sky130_fd_pr__special_nfet_latch ad=0.45 pd=2.8 as=0.189 ps=1.32 w=0.9 l=0.3
X1 a_n90_n42# a_n144_n130# a_n90_n244# w_n144_n252# sky130_fd_bs_flash__special_sonosfet_star ad=0.189 pd=1.32 as=0.513 ps=2.94 w=0.9 l=0.44
.ends

.subckt sonos_cell_mirrored sonos_cell_0/a_n144_n130# sonos_cell_0/a_n144_42# sonos_cell_1/dw_n144_n252#
+ w_160_160# sonos_cell_1/a_n144_42# sonos_cell_0/li_n144_n60# sonos_cell_1/a_n144_n130#
+ sonos_cell_1/a_n90_102# sonos_cell_1/a_n90_n244# sonos_cell_1/li_n144_n60#
Xsonos_cell_0 w_160_160# sonos_cell_0/a_n144_n130# sonos_cell_1/dw_n144_n252# sonos_cell_1/a_n90_n244#
+ sonos_cell_1/a_n90_102# sonos_cell_0/li_n144_n60# sonos_cell_0/a_n144_42# sonos_cell
Xsonos_cell_1 w_160_160# sonos_cell_1/a_n144_n130# sonos_cell_1/dw_n144_n252# sonos_cell_1/a_n90_n244#
+ sonos_cell_1/a_n90_102# sonos_cell_1/li_n144_n60# sonos_cell_1/a_n144_42# sonos_cell
.ends

.subckt sonos_8x8 w_n80_n96# dw_n80_n96#
Xsonos_cell_mirrored_0[0|0] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|0] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|0] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|0] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|1] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|1] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|1] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|1] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|2] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|2] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|2] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|2] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|3] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|3] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|3] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|3] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|4] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|4] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|4] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|4] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|5] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|5] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|5] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|5] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|6] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|6] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|6] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|6] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|7] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|7] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|7] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|7] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
.ends

.subckt sonos_array_50x50x64 w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96#
Xsonos_8x8_0[0|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
.ends

.subckt sonos_endcap_tb dw_n408_n1786# m1_n300_n1886# w_n120_n1786# w_n408_n1360#
+ a_n408_n922# a_n354_n1046#
X0 a_n354_n1046# a_n408_n922# a_n354_n1046# w_n408_n1360# sky130_fd_pr__nfet_01v8 ad=1.01 pd=5.84 as=0.45 ps=2.8 w=0.9 l=0.3
.ends

.subckt sonos_array_orig w_n498_n930#
Xsonos_endcap_tb_1[0] dw_0_n64# sonos_cell_2[3|0]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|0]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[1] dw_0_n64# sonos_cell_2[3|1]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|1]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[2] dw_0_n64# sonos_cell_2[3|2]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|2]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[3] dw_0_n64# sonos_cell_2[3|3]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|3]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[4] dw_0_n64# sonos_cell_2[3|4]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|4]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[5] dw_0_n64# sonos_cell_2[3|5]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|5]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[6] dw_0_n64# sonos_cell_2[3|6]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|6]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_1[7] dw_0_n64# sonos_cell_2[3|7]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_3/a_n72_n552# sonos_cell_2[3|7]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[0] dw_0_n64# sonos_cell_2[3|0]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|0]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[1] dw_0_n64# sonos_cell_2[3|1]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|1]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[2] dw_0_n64# sonos_cell_2[3|2]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|2]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[3] dw_0_n64# sonos_cell_2[3|3]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|3]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[4] dw_0_n64# sonos_cell_2[3|4]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|4]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[5] dw_0_n64# sonos_cell_2[3|5]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|5]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[6] dw_0_n64# sonos_cell_2[3|6]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|6]/a_n90_102# sonos_endcap_tb
Xsonos_endcap_tb_2[7] dw_0_n64# sonos_cell_2[3|7]/a_n90_n244# w_n498_n930# w_n498_n930#
+ sonos_array_corner_4/a_n72_n552# sonos_cell_2[3|7]/a_n90_102# sonos_endcap_tb
Xsonos_cell_1[0|0] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244# sonos_cell_2[3|0]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|0] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|0] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|0] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|1] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244# sonos_cell_2[3|1]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|1] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|1] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|1] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|2] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244# sonos_cell_2[3|2]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|2] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|2] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|2] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|3] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244# sonos_cell_2[3|3]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|3] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|3] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|3] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|4] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244# sonos_cell_2[3|4]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|4] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|4] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|4] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|5] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244# sonos_cell_2[3|5]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|5] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|5] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|5] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|6] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244# sonos_cell_2[3|6]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|6] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|6] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|6] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[0|7] w_n498_n930# a_0_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244# sonos_cell_2[3|7]/a_n90_102#
+ sonos_cell_1[0|7]/li_n144_n60# a_0_200# sonos_cell
Xsonos_cell_1[1|7] w_n498_n930# sonos_endcap_lr_1[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_1[1|7]/li_n144_n60# sonos_cell_1[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[2|7] w_n498_n930# sonos_endcap_lr_1[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_1[2|7]/li_n144_n60# sonos_cell_1[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_1[3|7] w_n498_n930# sonos_endcap_lr_1[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_1[3|7]/li_n144_n60# sonos_cell_1[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|0] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|0] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|0] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|0] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|0]/a_n90_n244#
+ sonos_cell_2[3|0]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|1] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|1] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|1] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|1] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|1]/a_n90_n244#
+ sonos_cell_2[3|1]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|2] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|2] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|2] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|2] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|2]/a_n90_n244#
+ sonos_cell_2[3|2]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|3] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|3] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|3] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|3] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|3]/a_n90_n244#
+ sonos_cell_2[3|3]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|4] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|4] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|4] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|4] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|4]/a_n90_n244#
+ sonos_cell_2[3|4]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|5] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|5] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|5] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|5] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|5]/a_n90_n244#
+ sonos_cell_2[3|5]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|6] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|6] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|6] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|6] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|6]/a_n90_n244#
+ sonos_cell_2[3|6]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[0|7] w_n498_n930# sonos_endcap_lr_2[3]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_2[0|7]/li_n144_n60# sonos_cell_2[0|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[1|7] w_n498_n930# sonos_endcap_lr_2[2]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_2[1|7]/li_n144_n60# sonos_cell_2[1|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[2|7] w_n498_n930# sonos_endcap_lr_2[1]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_2[2|7]/li_n144_n60# sonos_cell_2[2|7]/a_n144_42#
+ sonos_cell
Xsonos_cell_2[3|7] w_n498_n930# sonos_endcap_lr_2[0]/a_n72_28# dw_0_n64# sonos_cell_2[3|7]/a_n90_n244#
+ sonos_cell_2[3|7]/a_n90_102# sonos_cell_2[3|7]/li_n144_n60# sonos_cell_2[3|7]/a_n144_42#
+ sonos_cell
.ends

.subckt sonos_array_labeled VPB
Xsonos_array_orig_0 VPB sonos_array_orig
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xsonos_array_50x50x64_0 w_21434_30636# dw_21184_30386# sonos_array_50x50x64
Xsonos_array_labeled_0[0|0] sonos_array_labeled_0[0|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|0] sonos_array_labeled_0[1|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|0] sonos_array_labeled_0[2|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|0] sonos_array_labeled_0[3|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|0] sonos_array_labeled_0[4|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|0] sonos_array_labeled_0[5|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|0] sonos_array_labeled_0[6|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|0] sonos_array_labeled_0[7|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|0] sonos_array_labeled_0[8|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|0] sonos_array_labeled_0[9|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|0] sonos_array_labeled_0[10|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|0] sonos_array_labeled_0[11|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|0] sonos_array_labeled_0[12|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|0] sonos_array_labeled_0[13|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|0] sonos_array_labeled_0[14|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|0] sonos_array_labeled_0[15|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|0] sonos_array_labeled_0[16|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|0] sonos_array_labeled_0[17|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|0] sonos_array_labeled_0[18|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|0] sonos_array_labeled_0[19|0]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|1] sonos_array_labeled_0[0|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|1] sonos_array_labeled_0[1|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|1] sonos_array_labeled_0[2|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|1] sonos_array_labeled_0[3|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|1] sonos_array_labeled_0[4|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|1] sonos_array_labeled_0[5|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|1] sonos_array_labeled_0[6|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|1] sonos_array_labeled_0[7|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|1] sonos_array_labeled_0[8|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|1] sonos_array_labeled_0[9|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|1] sonos_array_labeled_0[10|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|1] sonos_array_labeled_0[11|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|1] sonos_array_labeled_0[12|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|1] sonos_array_labeled_0[13|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|1] sonos_array_labeled_0[14|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|1] sonos_array_labeled_0[15|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|1] sonos_array_labeled_0[16|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|1] sonos_array_labeled_0[17|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|1] sonos_array_labeled_0[18|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|1] sonos_array_labeled_0[19|1]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|2] sonos_array_labeled_0[0|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|2] sonos_array_labeled_0[1|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|2] sonos_array_labeled_0[2|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|2] sonos_array_labeled_0[3|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|2] sonos_array_labeled_0[4|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|2] sonos_array_labeled_0[5|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|2] sonos_array_labeled_0[6|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|2] sonos_array_labeled_0[7|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|2] sonos_array_labeled_0[8|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|2] sonos_array_labeled_0[9|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|2] sonos_array_labeled_0[10|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|2] sonos_array_labeled_0[11|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|2] sonos_array_labeled_0[12|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|2] sonos_array_labeled_0[13|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|2] sonos_array_labeled_0[14|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|2] sonos_array_labeled_0[15|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|2] sonos_array_labeled_0[16|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|2] sonos_array_labeled_0[17|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|2] sonos_array_labeled_0[18|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|2] sonos_array_labeled_0[19|2]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|3] sonos_array_labeled_0[0|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|3] sonos_array_labeled_0[1|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|3] sonos_array_labeled_0[2|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|3] sonos_array_labeled_0[3|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|3] sonos_array_labeled_0[4|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|3] sonos_array_labeled_0[5|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|3] sonos_array_labeled_0[6|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|3] sonos_array_labeled_0[7|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|3] sonos_array_labeled_0[8|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|3] sonos_array_labeled_0[9|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|3] sonos_array_labeled_0[10|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|3] sonos_array_labeled_0[11|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|3] sonos_array_labeled_0[12|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|3] sonos_array_labeled_0[13|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|3] sonos_array_labeled_0[14|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|3] sonos_array_labeled_0[15|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|3] sonos_array_labeled_0[16|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|3] sonos_array_labeled_0[17|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|3] sonos_array_labeled_0[18|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|3] sonos_array_labeled_0[19|3]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|4] sonos_array_labeled_0[0|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|4] sonos_array_labeled_0[1|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|4] sonos_array_labeled_0[2|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|4] sonos_array_labeled_0[3|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|4] sonos_array_labeled_0[4|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|4] sonos_array_labeled_0[5|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|4] sonos_array_labeled_0[6|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|4] sonos_array_labeled_0[7|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|4] sonos_array_labeled_0[8|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|4] sonos_array_labeled_0[9|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|4] sonos_array_labeled_0[10|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|4] sonos_array_labeled_0[11|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|4] sonos_array_labeled_0[12|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|4] sonos_array_labeled_0[13|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|4] sonos_array_labeled_0[14|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|4] sonos_array_labeled_0[15|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|4] sonos_array_labeled_0[16|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|4] sonos_array_labeled_0[17|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|4] sonos_array_labeled_0[18|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|4] sonos_array_labeled_0[19|4]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|5] sonos_array_labeled_0[0|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|5] sonos_array_labeled_0[1|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|5] sonos_array_labeled_0[2|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|5] sonos_array_labeled_0[3|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|5] sonos_array_labeled_0[4|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|5] sonos_array_labeled_0[5|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|5] sonos_array_labeled_0[6|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|5] sonos_array_labeled_0[7|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|5] sonos_array_labeled_0[8|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|5] sonos_array_labeled_0[9|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|5] sonos_array_labeled_0[10|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|5] sonos_array_labeled_0[11|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|5] sonos_array_labeled_0[12|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|5] sonos_array_labeled_0[13|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|5] sonos_array_labeled_0[14|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|5] sonos_array_labeled_0[15|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|5] sonos_array_labeled_0[16|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|5] sonos_array_labeled_0[17|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|5] sonos_array_labeled_0[18|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|5] sonos_array_labeled_0[19|5]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|6] sonos_array_labeled_0[0|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|6] sonos_array_labeled_0[1|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|6] sonos_array_labeled_0[2|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|6] sonos_array_labeled_0[3|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|6] sonos_array_labeled_0[4|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|6] sonos_array_labeled_0[5|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|6] sonos_array_labeled_0[6|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|6] sonos_array_labeled_0[7|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|6] sonos_array_labeled_0[8|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|6] sonos_array_labeled_0[9|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|6] sonos_array_labeled_0[10|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|6] sonos_array_labeled_0[11|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|6] sonos_array_labeled_0[12|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|6] sonos_array_labeled_0[13|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|6] sonos_array_labeled_0[14|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|6] sonos_array_labeled_0[15|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|6] sonos_array_labeled_0[16|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|6] sonos_array_labeled_0[17|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|6] sonos_array_labeled_0[18|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|6] sonos_array_labeled_0[19|6]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|7] sonos_array_labeled_0[0|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|7] sonos_array_labeled_0[1|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|7] sonos_array_labeled_0[2|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|7] sonos_array_labeled_0[3|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|7] sonos_array_labeled_0[4|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|7] sonos_array_labeled_0[5|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|7] sonos_array_labeled_0[6|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|7] sonos_array_labeled_0[7|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|7] sonos_array_labeled_0[8|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|7] sonos_array_labeled_0[9|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|7] sonos_array_labeled_0[10|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|7] sonos_array_labeled_0[11|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|7] sonos_array_labeled_0[12|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|7] sonos_array_labeled_0[13|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|7] sonos_array_labeled_0[14|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|7] sonos_array_labeled_0[15|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|7] sonos_array_labeled_0[16|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|7] sonos_array_labeled_0[17|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|7] sonos_array_labeled_0[18|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|7] sonos_array_labeled_0[19|7]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|8] sonos_array_labeled_0[0|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|8] sonos_array_labeled_0[1|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|8] sonos_array_labeled_0[2|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|8] sonos_array_labeled_0[3|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|8] sonos_array_labeled_0[4|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|8] sonos_array_labeled_0[5|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|8] sonos_array_labeled_0[6|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|8] sonos_array_labeled_0[7|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|8] sonos_array_labeled_0[8|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|8] sonos_array_labeled_0[9|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|8] sonos_array_labeled_0[10|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|8] sonos_array_labeled_0[11|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|8] sonos_array_labeled_0[12|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|8] sonos_array_labeled_0[13|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|8] sonos_array_labeled_0[14|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|8] sonos_array_labeled_0[15|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|8] sonos_array_labeled_0[16|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|8] sonos_array_labeled_0[17|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|8] sonos_array_labeled_0[18|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|8] sonos_array_labeled_0[19|8]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|9] sonos_array_labeled_0[0|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|9] sonos_array_labeled_0[1|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|9] sonos_array_labeled_0[2|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|9] sonos_array_labeled_0[3|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|9] sonos_array_labeled_0[4|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|9] sonos_array_labeled_0[5|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|9] sonos_array_labeled_0[6|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|9] sonos_array_labeled_0[7|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|9] sonos_array_labeled_0[8|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|9] sonos_array_labeled_0[9|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|9] sonos_array_labeled_0[10|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|9] sonos_array_labeled_0[11|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|9] sonos_array_labeled_0[12|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|9] sonos_array_labeled_0[13|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|9] sonos_array_labeled_0[14|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|9] sonos_array_labeled_0[15|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|9] sonos_array_labeled_0[16|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|9] sonos_array_labeled_0[17|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|9] sonos_array_labeled_0[18|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|9] sonos_array_labeled_0[19|9]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|10] sonos_array_labeled_0[0|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|10] sonos_array_labeled_0[1|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|10] sonos_array_labeled_0[2|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|10] sonos_array_labeled_0[3|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|10] sonos_array_labeled_0[4|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|10] sonos_array_labeled_0[5|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|10] sonos_array_labeled_0[6|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|10] sonos_array_labeled_0[7|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|10] sonos_array_labeled_0[8|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|10] sonos_array_labeled_0[9|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|10] sonos_array_labeled_0[10|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|10] sonos_array_labeled_0[11|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|10] sonos_array_labeled_0[12|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|10] sonos_array_labeled_0[13|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|10] sonos_array_labeled_0[14|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|10] sonos_array_labeled_0[15|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|10] sonos_array_labeled_0[16|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|10] sonos_array_labeled_0[17|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|10] sonos_array_labeled_0[18|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|10] sonos_array_labeled_0[19|10]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|11] sonos_array_labeled_0[0|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|11] sonos_array_labeled_0[1|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|11] sonos_array_labeled_0[2|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|11] sonos_array_labeled_0[3|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|11] sonos_array_labeled_0[4|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|11] sonos_array_labeled_0[5|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|11] sonos_array_labeled_0[6|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|11] sonos_array_labeled_0[7|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|11] sonos_array_labeled_0[8|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|11] sonos_array_labeled_0[9|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|11] sonos_array_labeled_0[10|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|11] sonos_array_labeled_0[11|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|11] sonos_array_labeled_0[12|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|11] sonos_array_labeled_0[13|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|11] sonos_array_labeled_0[14|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|11] sonos_array_labeled_0[15|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|11] sonos_array_labeled_0[16|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|11] sonos_array_labeled_0[17|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|11] sonos_array_labeled_0[18|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|11] sonos_array_labeled_0[19|11]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|12] sonos_array_labeled_0[0|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|12] sonos_array_labeled_0[1|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|12] sonos_array_labeled_0[2|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|12] sonos_array_labeled_0[3|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|12] sonos_array_labeled_0[4|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|12] sonos_array_labeled_0[5|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|12] sonos_array_labeled_0[6|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|12] sonos_array_labeled_0[7|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|12] sonos_array_labeled_0[8|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|12] sonos_array_labeled_0[9|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|12] sonos_array_labeled_0[10|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|12] sonos_array_labeled_0[11|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|12] sonos_array_labeled_0[12|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|12] sonos_array_labeled_0[13|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|12] sonos_array_labeled_0[14|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|12] sonos_array_labeled_0[15|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|12] sonos_array_labeled_0[16|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|12] sonos_array_labeled_0[17|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|12] sonos_array_labeled_0[18|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|12] sonos_array_labeled_0[19|12]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|13] sonos_array_labeled_0[0|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|13] sonos_array_labeled_0[1|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|13] sonos_array_labeled_0[2|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|13] sonos_array_labeled_0[3|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|13] sonos_array_labeled_0[4|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|13] sonos_array_labeled_0[5|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|13] sonos_array_labeled_0[6|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|13] sonos_array_labeled_0[7|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|13] sonos_array_labeled_0[8|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|13] sonos_array_labeled_0[9|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|13] sonos_array_labeled_0[10|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|13] sonos_array_labeled_0[11|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|13] sonos_array_labeled_0[12|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|13] sonos_array_labeled_0[13|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|13] sonos_array_labeled_0[14|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|13] sonos_array_labeled_0[15|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|13] sonos_array_labeled_0[16|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|13] sonos_array_labeled_0[17|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|13] sonos_array_labeled_0[18|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|13] sonos_array_labeled_0[19|13]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|14] sonos_array_labeled_0[0|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|14] sonos_array_labeled_0[1|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|14] sonos_array_labeled_0[2|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|14] sonos_array_labeled_0[3|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|14] sonos_array_labeled_0[4|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|14] sonos_array_labeled_0[5|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|14] sonos_array_labeled_0[6|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|14] sonos_array_labeled_0[7|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|14] sonos_array_labeled_0[8|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|14] sonos_array_labeled_0[9|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|14] sonos_array_labeled_0[10|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|14] sonos_array_labeled_0[11|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|14] sonos_array_labeled_0[12|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|14] sonos_array_labeled_0[13|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|14] sonos_array_labeled_0[14|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|14] sonos_array_labeled_0[15|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|14] sonos_array_labeled_0[16|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|14] sonos_array_labeled_0[17|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|14] sonos_array_labeled_0[18|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|14] sonos_array_labeled_0[19|14]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|15] sonos_array_labeled_0[0|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|15] sonos_array_labeled_0[1|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|15] sonos_array_labeled_0[2|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|15] sonos_array_labeled_0[3|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|15] sonos_array_labeled_0[4|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|15] sonos_array_labeled_0[5|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|15] sonos_array_labeled_0[6|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|15] sonos_array_labeled_0[7|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|15] sonos_array_labeled_0[8|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|15] sonos_array_labeled_0[9|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|15] sonos_array_labeled_0[10|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|15] sonos_array_labeled_0[11|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|15] sonos_array_labeled_0[12|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|15] sonos_array_labeled_0[13|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|15] sonos_array_labeled_0[14|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|15] sonos_array_labeled_0[15|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|15] sonos_array_labeled_0[16|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|15] sonos_array_labeled_0[17|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|15] sonos_array_labeled_0[18|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|15] sonos_array_labeled_0[19|15]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|16] sonos_array_labeled_0[0|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|16] sonos_array_labeled_0[1|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|16] sonos_array_labeled_0[2|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|16] sonos_array_labeled_0[3|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|16] sonos_array_labeled_0[4|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|16] sonos_array_labeled_0[5|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|16] sonos_array_labeled_0[6|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|16] sonos_array_labeled_0[7|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|16] sonos_array_labeled_0[8|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|16] sonos_array_labeled_0[9|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|16] sonos_array_labeled_0[10|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|16] sonos_array_labeled_0[11|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|16] sonos_array_labeled_0[12|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|16] sonos_array_labeled_0[13|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|16] sonos_array_labeled_0[14|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|16] sonos_array_labeled_0[15|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|16] sonos_array_labeled_0[16|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|16] sonos_array_labeled_0[17|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|16] sonos_array_labeled_0[18|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|16] sonos_array_labeled_0[19|16]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|17] sonos_array_labeled_0[0|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|17] sonos_array_labeled_0[1|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|17] sonos_array_labeled_0[2|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|17] sonos_array_labeled_0[3|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|17] sonos_array_labeled_0[4|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|17] sonos_array_labeled_0[5|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|17] sonos_array_labeled_0[6|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|17] sonos_array_labeled_0[7|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|17] sonos_array_labeled_0[8|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|17] sonos_array_labeled_0[9|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|17] sonos_array_labeled_0[10|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|17] sonos_array_labeled_0[11|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|17] sonos_array_labeled_0[12|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|17] sonos_array_labeled_0[13|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|17] sonos_array_labeled_0[14|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|17] sonos_array_labeled_0[15|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|17] sonos_array_labeled_0[16|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|17] sonos_array_labeled_0[17|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|17] sonos_array_labeled_0[18|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|17] sonos_array_labeled_0[19|17]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|18] sonos_array_labeled_0[0|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|18] sonos_array_labeled_0[1|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|18] sonos_array_labeled_0[2|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|18] sonos_array_labeled_0[3|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|18] sonos_array_labeled_0[4|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|18] sonos_array_labeled_0[5|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|18] sonos_array_labeled_0[6|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|18] sonos_array_labeled_0[7|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|18] sonos_array_labeled_0[8|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|18] sonos_array_labeled_0[9|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|18] sonos_array_labeled_0[10|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|18] sonos_array_labeled_0[11|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|18] sonos_array_labeled_0[12|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|18] sonos_array_labeled_0[13|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|18] sonos_array_labeled_0[14|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|18] sonos_array_labeled_0[15|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|18] sonos_array_labeled_0[16|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|18] sonos_array_labeled_0[17|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|18] sonos_array_labeled_0[18|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|18] sonos_array_labeled_0[19|18]/VPB sonos_array_labeled
Xsonos_array_labeled_0[0|19] sonos_array_labeled_0[0|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[1|19] sonos_array_labeled_0[1|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[2|19] sonos_array_labeled_0[2|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[3|19] sonos_array_labeled_0[3|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[4|19] sonos_array_labeled_0[4|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[5|19] sonos_array_labeled_0[5|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[6|19] sonos_array_labeled_0[6|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[7|19] sonos_array_labeled_0[7|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[8|19] sonos_array_labeled_0[8|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[9|19] sonos_array_labeled_0[9|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[10|19] sonos_array_labeled_0[10|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[11|19] sonos_array_labeled_0[11|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[12|19] sonos_array_labeled_0[12|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[13|19] sonos_array_labeled_0[13|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[14|19] sonos_array_labeled_0[14|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[15|19] sonos_array_labeled_0[15|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[16|19] sonos_array_labeled_0[16|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[17|19] sonos_array_labeled_0[17|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[18|19] sonos_array_labeled_0[18|19]/VPB sonos_array_labeled
Xsonos_array_labeled_0[19|19] sonos_array_labeled_0[19|19]/VPB sonos_array_labeled
.ends

