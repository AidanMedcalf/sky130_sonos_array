magic
tech sky130A
timestamp 1685134277
<< metal3 >>
rect -25 16 25 24
rect -25 -16 -16 16
rect 16 -16 25 16
rect -25 -24 25 -16
<< via3 >>
rect -16 -16 16 16
<< via4 >>
rect -59 16 59 59
rect -59 -16 -16 16
rect -16 -16 16 16
rect 16 -16 59 16
rect -59 -59 59 -16
<< metal5 >>
rect -100 59 100 100
rect -100 -59 -59 59
rect 59 -59 100 59
rect -100 -100 100 -59
<< glass >>
rect -90 -90 90 90
<< end >>
