magic
tech sky130A
magscale 1 2
timestamp 1663459791
<< error_p >>
rect 352 485 520 941
rect 358 429 404 441
rect 468 429 514 441
rect 358 395 364 429
rect 468 395 474 429
rect 358 383 404 395
rect 468 383 514 395
rect 520 341 952 485
use sky130_fd_bs_flash__special_sonosfet_star_8ZR9Z2  sky130_fd_bs_flash__special_sonosfet_star_8ZR9Z2_0
timestamp 1663459791
transform 1 0 436 0 1 411
box -84 -70 516 530
<< end >>
