magic
tech sky130A
timestamp 1686079789
<< dnwell >>
rect -40 -48 1210 1490
use sonos_8x8  sonos_8x8_0
timestamp 1686079789
transform 1 0 0 0 1 0
box -40 -48 1308 1490
<< end >>
