magic
tech sky130A
magscale 1 2
timestamp 1663459876
<< error_p >>
rect 0 1152 938 1608
rect 0 144 1370 1152
rect 6 88 52 100
rect 116 88 162 100
rect 6 54 12 88
rect 116 54 122 88
rect 6 42 52 54
rect 116 42 162 54
rect 168 0 1370 144
use sonos_small  sonos_small_0
array 0 7 110 0 7 144
timestamp 1663459791
transform 1 0 -352 0 1 -341
box 352 341 952 941
<< end >>
