* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_bs_flash__special_sonosfet_star w_n436_n442# a_n33_36# dw_n436_n442#
+ a_22_n76# a_n84_n76#
X0 a_22_n76# a_n33_36# a_n84_n76# w_n436_n442# sky130_fd_bs_flash__special_sonosfet_star ad=1.395e+11p pd=1.52e+06u as=1.395e+11p ps=1.52e+06u w=450000u l=220000u
.ends

.subckt sonos_cell w_n144_n252# a_n144_n130# dw_n144_n252# a_n90_n244# a_n90_102#
+ li_n144_n60# a_n144_42#
X0 a_n90_102# a_n144_42# a_n90_n42# w_n144_n252# sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=3.78e+11p ps=2.64e+06u w=900000u l=300000u
X1 a_n90_n42# a_n144_n130# a_n90_n244# w_n144_n252# sky130_fd_bs_flash__special_sonosfet_star ad=0p pd=0u as=5.13e+11p ps=2.94e+06u w=900000u l=440000u
.ends

.subckt sonos_cell_mirrored sonos_cell_0/a_n144_n130# sonos_cell_0/a_n144_42# sonos_cell_1/dw_n144_n252#
+ w_160_160# sonos_cell_1/a_n144_42# sonos_cell_0/li_n144_n60# sonos_cell_1/a_n144_n130#
+ sonos_cell_1/a_n90_102# sonos_cell_1/a_n90_n244# sonos_cell_1/li_n144_n60#
Xsonos_cell_0 w_160_160# sonos_cell_0/a_n144_n130# sonos_cell_1/dw_n144_n252# sonos_cell_1/a_n90_n244#
+ sonos_cell_1/a_n90_102# sonos_cell_0/li_n144_n60# sonos_cell_0/a_n144_42# sonos_cell
Xsonos_cell_1 w_160_160# sonos_cell_1/a_n144_n130# sonos_cell_1/dw_n144_n252# sonos_cell_1/a_n90_n244#
+ sonos_cell_1/a_n90_102# sonos_cell_1/li_n144_n60# sonos_cell_1/a_n144_42# sonos_cell
.ends

.subckt sonos_8x8 w_n80_n96# dw_n80_n96#
Xsonos_cell_mirrored_0[0|0] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|0] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|0] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|0] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|1] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|1] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|1] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|1] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|2] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|2] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|2] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|2] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|3] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|3] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|3] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|3] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|4] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|4] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|4] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|4] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|5] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|5] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|5] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|5] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|6] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|6] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|6] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|6] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[0|7] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[1|7] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[2|7] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
Xsonos_cell_mirrored_0[3|7] w_n80_n96# w_n80_n96# dw_n80_n96# w_n80_n96# w_n80_n96#
+ w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# w_n80_n96# sonos_cell_mirrored
.ends

.subckt sonos_array_240x250x64 w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96#
Xsonos_8x8_0[0|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|0] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|1] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|2] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|3] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|4] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|5] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|6] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|7] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|8] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|9] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|10] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|11] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|12] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|13] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|14] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|15] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|16] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|17] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|18] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|19] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|20] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|21] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|22] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|23] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|24] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|25] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|26] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|27] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|28] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|29] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|30] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|31] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|32] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|33] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|34] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|35] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|36] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|37] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|38] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|39] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|40] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|41] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|42] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|43] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|44] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|45] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|46] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|47] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|48] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|49] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|50] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|51] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|52] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|53] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|54] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|55] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|56] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|57] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|58] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|59] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|60] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|61] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|62] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|63] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|64] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|65] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|66] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|67] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|68] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|69] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|70] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|71] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|72] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|73] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|74] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|75] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|76] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|77] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|78] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|79] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|80] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|81] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|82] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|83] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|84] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|85] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|86] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|87] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|88] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|89] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|90] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|91] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|92] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|93] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|94] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|95] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|96] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|97] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|98] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|99] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|100] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|101] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|102] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|103] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|104] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|105] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|106] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|107] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|108] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|109] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|110] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|111] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|112] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|113] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|114] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|115] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|116] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|117] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|118] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|119] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|120] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|121] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|122] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|123] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|124] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|125] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|126] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|127] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|128] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|129] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|130] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|131] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|132] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|133] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|134] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|135] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|136] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|137] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|138] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|139] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|140] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|141] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|142] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|143] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|144] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|145] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|146] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|147] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|148] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|149] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|150] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|151] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|152] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|153] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|154] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|155] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|156] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|157] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|158] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|159] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|160] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|161] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|162] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|163] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|164] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|165] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|166] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|167] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|168] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|169] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|170] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|171] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|172] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|173] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|174] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|175] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|176] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|177] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|178] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|179] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|180] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|181] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|182] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|183] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|184] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|185] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|186] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|187] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|188] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|189] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|190] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|191] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|192] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|193] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|194] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|195] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|196] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|197] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|198] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|199] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|200] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|201] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|202] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|203] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|204] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|205] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|206] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|207] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|208] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|209] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|210] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|211] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|212] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|213] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|214] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|215] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|216] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|217] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|218] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|219] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|220] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|221] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|222] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|223] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|224] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|225] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|226] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|227] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|228] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|229] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|230] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|231] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|232] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|233] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[0|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[1|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[2|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[3|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[4|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[5|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[6|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[7|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[8|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[9|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[10|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[11|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[12|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[13|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[14|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[15|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[16|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[17|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[18|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[19|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[20|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[21|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[22|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[23|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[24|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[25|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[26|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[27|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[28|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[29|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[30|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[31|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[32|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[33|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[34|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[35|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[36|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[37|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[38|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[39|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[40|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[41|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[42|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[43|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[44|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[45|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[46|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[47|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[48|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[49|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[50|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[51|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[52|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[53|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[54|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[55|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[56|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[57|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[58|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[59|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[60|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[61|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[62|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[63|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[64|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[65|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[66|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[67|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[68|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[69|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[70|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[71|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[72|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[73|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[74|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[75|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[76|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[77|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[78|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[79|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[80|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[81|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[82|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[83|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[84|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[85|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[86|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[87|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[88|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[89|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[90|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[91|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[92|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[93|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[94|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[95|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[96|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[97|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[98|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[99|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[100|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[101|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[102|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[103|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[104|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[105|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[106|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[107|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[108|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[109|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[110|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[111|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[112|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[113|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[114|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[115|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[116|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[117|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[118|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[119|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[120|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[121|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[122|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[123|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[124|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[125|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[126|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[127|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[128|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[129|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[130|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[131|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[132|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[133|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[134|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[135|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[136|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[137|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[138|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[139|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[140|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[141|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[142|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[143|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[144|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[145|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[146|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[147|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[148|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[149|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[150|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[151|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[152|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[153|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[154|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[155|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[156|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[157|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[158|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[159|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[160|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[161|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[162|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[163|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[164|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[165|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[166|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[167|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[168|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[169|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[170|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[171|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[172|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[173|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[174|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[175|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[176|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[177|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[178|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[179|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[180|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[181|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[182|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[183|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[184|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[185|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[186|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[187|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[188|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[189|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[190|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[191|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[192|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[193|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[194|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[195|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[196|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[197|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[198|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[199|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[200|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[201|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[202|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[203|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[204|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[205|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[206|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[207|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[208|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[209|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[210|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[211|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[212|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[213|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
Xsonos_8x8_0[214|234] w_n80_n96# sonos_8x8_0[9|9]/dw_n80_n96# sonos_8x8
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xsky130_fd_bs_flash__special_sonosfet_star_0 vssa1 io_analog[9] vdda1 io_analog[8]
+ io_analog[10] sky130_fd_bs_flash__special_sonosfet_star
Xsky130_fd_bs_flash__special_sonosfet_star_1 io_analog[7] io_analog[5] vdda1 io_analog[4]
+ io_analog[6] sky130_fd_bs_flash__special_sonosfet_star
Xsky130_fd_bs_flash__special_sonosfet_star_2 io_analog[3] io_analog[1] vdda1 io_analog[0]
+ io_analog[2] sky130_fd_bs_flash__special_sonosfet_star
Xsonos_array_240x250x64_0 vssa2 vdda2 sonos_array_240x250x64
.ends

