magic
tech sky130A
timestamp 1663486910
use sonos_8x8  sonos_8x8_0
array 0 234 1225 0 214 1513
timestamp 1663485803
transform 1 0 0 0 1 0
box -40 -48 1308 1490
<< end >>
