magic
tech sky130A
timestamp 1663450679
<< error_s >>
rect -152 1461 1337 1604
rect -152 -19 -9 1461
rect 27 1337 117 1381
rect 171 1337 261 1381
rect 315 1337 405 1381
rect 459 1337 549 1381
rect 603 1337 693 1381
rect 747 1337 837 1381
rect 891 1337 981 1381
rect 1035 1337 1125 1381
rect 27 1099 117 1143
rect 171 1099 261 1143
rect 315 1099 405 1143
rect 459 1099 549 1143
rect 603 1099 693 1143
rect 747 1099 837 1143
rect 891 1099 981 1143
rect 1035 1099 1125 1143
rect 27 991 117 1035
rect 171 991 261 1035
rect 315 991 405 1035
rect 459 991 549 1035
rect 603 991 693 1035
rect 747 991 837 1035
rect 891 991 981 1035
rect 1035 991 1125 1035
rect 27 753 117 797
rect 171 753 261 797
rect 315 753 405 797
rect 459 753 549 797
rect 603 753 693 797
rect 747 753 837 797
rect 891 753 981 797
rect 1035 753 1125 797
rect 27 645 117 689
rect 171 645 261 689
rect 315 645 405 689
rect 459 645 549 689
rect 603 645 693 689
rect 747 645 837 689
rect 891 645 981 689
rect 1035 645 1125 689
rect 27 407 117 451
rect 171 407 261 451
rect 315 407 405 451
rect 459 407 549 451
rect 603 407 693 451
rect 747 407 837 451
rect 891 407 981 451
rect 1035 407 1125 451
rect 27 299 117 343
rect 171 299 261 343
rect 315 299 405 343
rect 459 299 549 343
rect 603 299 693 343
rect 747 299 837 343
rect 891 299 981 343
rect 1035 299 1125 343
rect 27 61 117 105
rect 171 61 261 105
rect 315 61 405 105
rect 459 61 549 105
rect 603 61 693 105
rect 747 61 837 105
rect 891 61 981 105
rect 1035 61 1125 105
rect 1194 -19 1337 1461
rect -152 -162 1337 -19
<< dnwell >>
rect -112 -122 1297 1564
<< psubdiff >>
rect -112 1515 0 1564
rect 1173 1515 1297 1564
rect -112 1442 -63 1515
rect 1248 1442 1297 1515
rect -112 -73 -63 0
rect 1248 -73 1297 0
rect -112 -122 0 -73
rect 1173 -122 1297 -73
<< locali >>
rect -100 1527 1285 1552
rect -100 -85 -75 1527
rect 1260 -85 1285 1527
rect -100 -110 1285 -85
use sonos_8x8  sonos_8x8_0
timestamp 1663450679
transform 1 0 0 0 1 0
box -40 -40 1308 1482
use sonos_cell_hshort  sonos_cell_hshort_0
array 0 0 300 0 3 346
timestamp 1663450679
transform 1 0 0 0 1 0
box -152 -40 188 444
use sonos_cell_hshort  sonos_cell_hshort_1
array 0 0 -300 0 3 346
timestamp 1663450679
transform -1 0 1185 0 1 0
box -152 -40 188 444
use sonos_cell_vshort  sonos_cell_vshort_0
array 0 7 144 0 0 58
timestamp 1663450679
transform 1 0 0 0 1 1038
box -40 359 300 699
use sonos_cell_vshort  sonos_cell_vshort_1
array 0 7 144 0 0 -58
timestamp 1663450679
transform 1 0 0 0 -1 404
box -40 359 300 699
<< end >>
