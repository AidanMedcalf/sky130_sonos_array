magic
tech sky130A
timestamp 1663485803
<< error_s >>
rect 224 80 380 484
use sonos_cell  sonos_cell_0
timestamp 1663485803
transform 1 0 152 0 1 206
box -72 -126 228 174
use sonos_cell  sonos_cell_1
timestamp 1663485803
transform 1 0 152 0 -1 358
box -72 -126 228 174
<< properties >>
string FIXED_BBOX 80 80 240 484
<< end >>
