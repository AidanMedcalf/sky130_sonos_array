magic
tech sky130A
timestamp 1686079789
<< error_p >>
rect -530 134 -449 152
rect -111 134 -36 145
rect -512 116 -467 134
rect -512 -212 -467 -194
rect -249 -212 0 134
rect -530 -230 -449 -212
<< dnwell >>
rect -462 -212 0 134
<< nwell >>
rect -548 -212 -249 134
<< srampvar >>
rect -111 100 -36 130
rect -111 14 -36 58
rect -111 -94 -36 -50
rect -111 -166 -36 -136
<< psubdiff >>
rect -111 130 -36 134
rect -111 58 -36 100
rect -111 -1 -36 14
rect -111 -35 -91 -1
rect -57 -35 -36 -1
rect -111 -50 -36 -35
rect -111 -136 -36 -94
rect -111 -173 -36 -166
rect -111 -207 -91 -173
rect -57 -207 -36 -173
rect -111 -212 -36 -207
<< nsubdiff >>
rect -512 121 -467 134
rect -512 -161 -507 121
rect -473 -161 -467 121
rect -512 -212 -467 -161
<< psubdiffcont >>
rect -91 -35 -57 -1
rect -91 -207 -57 -173
<< nsubdiffcont >>
rect -507 -161 -473 121
<< poly >>
rect -133 100 -111 130
rect -36 100 0 130
rect -308 64 -254 81
rect -308 30 -298 64
rect -264 58 -254 64
rect -264 30 -111 58
rect -308 14 -111 30
rect -36 14 0 58
rect -308 -50 -254 -34
rect -308 -51 -111 -50
rect -308 -85 -298 -51
rect -264 -85 -111 -51
rect -308 -94 -111 -85
rect -36 -94 0 -50
rect -308 -101 -254 -94
rect -227 -153 -111 -136
rect -227 -187 -217 -153
rect -183 -166 -111 -153
rect -36 -166 0 -136
rect -183 -187 -173 -166
rect -227 -203 -173 -187
<< polycont >>
rect -298 30 -264 64
rect -298 -85 -264 -51
rect -217 -187 -183 -153
<< locali >>
rect -507 121 -473 134
rect -298 64 -264 80
rect -298 14 -264 23
rect -210 66 0 83
rect -210 32 -199 66
rect -165 49 0 66
rect -165 32 -152 49
rect -210 19 -152 32
rect -91 -1 -57 15
rect -298 -51 -264 -35
rect -91 -51 -57 -35
rect -210 -72 -152 -55
rect -210 -106 -199 -72
rect -165 -85 -152 -72
rect -165 -106 0 -85
rect -210 -119 0 -106
rect -507 -212 -473 -161
rect -264 -187 -217 -153
rect -183 -187 -167 -153
rect -91 -173 -57 -157
rect -91 -223 -57 -207
<< viali >>
rect -298 30 -264 57
rect -298 23 -264 30
rect -199 32 -165 66
rect -91 -35 -57 -1
rect -298 -85 -264 -79
rect -298 -113 -264 -85
rect -199 -106 -165 -72
rect -298 -187 -264 -153
rect -91 -207 -57 -173
<< metal1 >>
rect -512 91 -177 125
rect -211 83 -177 91
rect -211 66 -152 83
rect -310 57 -252 63
rect -512 23 -298 57
rect -264 23 -252 57
rect -211 32 -199 66
rect -165 32 -152 66
rect -211 26 -152 32
rect -310 17 -252 23
rect -111 -1 -50 134
rect -512 -45 -177 -11
rect -210 -55 -177 -45
rect -111 -35 -91 -1
rect -57 -35 -50 -1
rect -210 -72 -152 -55
rect -310 -79 -252 -73
rect -512 -113 -298 -79
rect -264 -113 -252 -79
rect -310 -119 -252 -113
rect -210 -106 -199 -72
rect -165 -106 -152 -72
rect -210 -119 -152 -106
rect -310 -153 -252 -147
rect -512 -187 -298 -153
rect -264 -187 -252 -153
rect -310 -193 -252 -187
rect -111 -173 -50 -35
rect -111 -207 -91 -173
rect -57 -207 -50 -173
rect -111 -214 -50 -207
<< end >>
